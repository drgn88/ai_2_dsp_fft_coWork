`timescale 1ns / 1ps

module rom_twf_gen #(
    parameter ROM_DEPTH = 512,
    parameter TWF_WIDTH = 9,
    parameter ADDR_WIDTH = 9,
    parameter OFFSET = 64
) (
    // input clk,
    input [ADDR_WIDTH-1:0] addr,
    input en,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_R_add,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_Q_add,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_R_sub,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_Q_sub
);

    logic signed [TWF_WIDTH-1:0] rom_real_data[ROM_DEPTH-1:0];
    logic signed [TWF_WIDTH-1:0] rom_imag_data[ROM_DEPTH-1:0];

    always @(*) begin
            if(en) begin
            rom_real_data[0] = 128;
            rom_real_data[1] = 128;
            rom_real_data[2] = 128;
            rom_real_data[3] = 128;
            rom_real_data[4] = 128;
            rom_real_data[5] = 128;
            rom_real_data[6] = 128;
            rom_real_data[7] = 128;
            rom_real_data[8] = 128;
            rom_real_data[9] = 128;
            rom_real_data[10] = 128;
            rom_real_data[11] = 128;
            rom_real_data[12] = 128;
            rom_real_data[13] = 128;
            rom_real_data[14] = 128;
            rom_real_data[15] = 128;
            rom_real_data[16] = 128;
            rom_real_data[17] = 128;
            rom_real_data[18] = 128;
            rom_real_data[19] = 128;
            rom_real_data[20] = 128;
            rom_real_data[21] = 128;
            rom_real_data[22] = 128;
            rom_real_data[23] = 128;
            rom_real_data[24] = 128;
            rom_real_data[25] = 128;
            rom_real_data[26] = 128;
            rom_real_data[27] = 128;
            rom_real_data[28] = 128;
            rom_real_data[29] = 128;
            rom_real_data[30] = 128;
            rom_real_data[31] = 128;
            rom_real_data[32] = 128;
            rom_real_data[33] = 128;
            rom_real_data[34] = 128;
            rom_real_data[35] = 128;
            rom_real_data[36] = 128;
            rom_real_data[37] = 128;
            rom_real_data[38] = 128;
            rom_real_data[39] = 128;
            rom_real_data[40] = 128;
            rom_real_data[41] = 128;
            rom_real_data[42] = 128;
            rom_real_data[43] = 128;
            rom_real_data[44] = 128;
            rom_real_data[45] = 128;
            rom_real_data[46] = 128;
            rom_real_data[47] = 128;
            rom_real_data[48] = 128;
            rom_real_data[49] = 128;
            rom_real_data[50] = 128;
            rom_real_data[51] = 128;
            rom_real_data[52] = 128;
            rom_real_data[53] = 128;
            rom_real_data[54] = 128;
            rom_real_data[55] = 128;
            rom_real_data[56] = 128;
            rom_real_data[57] = 128;
            rom_real_data[58] = 128;
            rom_real_data[59] = 128;
            rom_real_data[60] = 128;
            rom_real_data[61] = 128;
            rom_real_data[62] = 128;
            rom_real_data[63] = 128;
            rom_real_data[64] = 128;
            rom_real_data[65] = 128;
            rom_real_data[66] = 127;
            rom_real_data[67] = 127;
            rom_real_data[68] = 126;
            rom_real_data[69] = 124;
            rom_real_data[70] = 122;
            rom_real_data[71] = 121;
            rom_real_data[72] = 118;
            rom_real_data[73] = 116;
            rom_real_data[74] = 113;
            rom_real_data[75] = 110;
            rom_real_data[76] = 106;
            rom_real_data[77] = 103;
            rom_real_data[78] = 99;
            rom_real_data[79] = 95;
            rom_real_data[80] = 91;
            rom_real_data[81] = 86;
            rom_real_data[82] = 81;
            rom_real_data[83] = 76;
            rom_real_data[84] = 71;
            rom_real_data[85] = 66;
            rom_real_data[86] = 60;
            rom_real_data[87] = 55;
            rom_real_data[88] = 49;
            rom_real_data[89] = 43;
            rom_real_data[90] = 37;
            rom_real_data[91] = 31;
            rom_real_data[92] = 25;
            rom_real_data[93] = 19;
            rom_real_data[94] = 13;
            rom_real_data[95] = 6;
            rom_real_data[96] = 0;
            rom_real_data[97] = -6;
            rom_real_data[98] = -13;
            rom_real_data[99] = -19;
            rom_real_data[100] = -25;
            rom_real_data[101] = -31;
            rom_real_data[102] = -37;
            rom_real_data[103] = -43;
            rom_real_data[104] = -49;
            rom_real_data[105] = -55;
            rom_real_data[106] = -60;
            rom_real_data[107] = -66;
            rom_real_data[108] = -71;
            rom_real_data[109] = -76;
            rom_real_data[110] = -81;
            rom_real_data[111] = -86;
            rom_real_data[112] = -91;
            rom_real_data[113] = -95;
            rom_real_data[114] = -99;
            rom_real_data[115] = -103;
            rom_real_data[116] = -106;
            rom_real_data[117] = -110;
            rom_real_data[118] = -113;
            rom_real_data[119] = -116;
            rom_real_data[120] = -118;
            rom_real_data[121] = -121;
            rom_real_data[122] = -122;
            rom_real_data[123] = -124;
            rom_real_data[124] = -126;
            rom_real_data[125] = -127;
            rom_real_data[126] = -127;
            rom_real_data[127] = -128;
            rom_real_data[128] = 128;
            rom_real_data[129] = 128;
            rom_real_data[130] = 128;
            rom_real_data[131] = 128;
            rom_real_data[132] = 127;
            rom_real_data[133] = 127;
            rom_real_data[134] = 127;
            rom_real_data[135] = 126;
            rom_real_data[136] = 126;
            rom_real_data[137] = 125;
            rom_real_data[138] = 124;
            rom_real_data[139] = 123;
            rom_real_data[140] = 122;
            rom_real_data[141] = 122;
            rom_real_data[142] = 121;
            rom_real_data[143] = 119;
            rom_real_data[144] = 118;
            rom_real_data[145] = 117;
            rom_real_data[146] = 116;
            rom_real_data[147] = 114;
            rom_real_data[148] = 113;
            rom_real_data[149] = 111;
            rom_real_data[150] = 110;
            rom_real_data[151] = 108;
            rom_real_data[152] = 106;
            rom_real_data[153] = 105;
            rom_real_data[154] = 103;
            rom_real_data[155] = 101;
            rom_real_data[156] = 99;
            rom_real_data[157] = 97;
            rom_real_data[158] = 95;
            rom_real_data[159] = 93;
            rom_real_data[160] = 91;
            rom_real_data[161] = 88;
            rom_real_data[162] = 86;
            rom_real_data[163] = 84;
            rom_real_data[164] = 81;
            rom_real_data[165] = 79;
            rom_real_data[166] = 76;
            rom_real_data[167] = 74;
            rom_real_data[168] = 71;
            rom_real_data[169] = 68;
            rom_real_data[170] = 66;
            rom_real_data[171] = 63;
            rom_real_data[172] = 60;
            rom_real_data[173] = 58;
            rom_real_data[174] = 55;
            rom_real_data[175] = 52;
            rom_real_data[176] = 49;
            rom_real_data[177] = 46;
            rom_real_data[178] = 43;
            rom_real_data[179] = 40;
            rom_real_data[180] = 37;
            rom_real_data[181] = 34;
            rom_real_data[182] = 31;
            rom_real_data[183] = 28;
            rom_real_data[184] = 25;
            rom_real_data[185] = 22;
            rom_real_data[186] = 19;
            rom_real_data[187] = 16;
            rom_real_data[188] = 13;
            rom_real_data[189] = 9;
            rom_real_data[190] = 6;
            rom_real_data[191] = 3;
            rom_real_data[192] = 128;
            rom_real_data[193] = 128;
            rom_real_data[194] = 127;
            rom_real_data[195] = 125;
            rom_real_data[196] = 122;
            rom_real_data[197] = 119;
            rom_real_data[198] = 116;
            rom_real_data[199] = 111;
            rom_real_data[200] = 106;
            rom_real_data[201] = 101;
            rom_real_data[202] = 95;
            rom_real_data[203] = 88;
            rom_real_data[204] = 81;
            rom_real_data[205] = 74;
            rom_real_data[206] = 66;
            rom_real_data[207] = 58;
            rom_real_data[208] = 49;
            rom_real_data[209] = 40;
            rom_real_data[210] = 31;
            rom_real_data[211] = 22;
            rom_real_data[212] = 13;
            rom_real_data[213] = 3;
            rom_real_data[214] = -6;
            rom_real_data[215] = -16;
            rom_real_data[216] = -25;
            rom_real_data[217] = -34;
            rom_real_data[218] = -43;
            rom_real_data[219] = -52;
            rom_real_data[220] = -60;
            rom_real_data[221] = -68;
            rom_real_data[222] = -76;
            rom_real_data[223] = -84;
            rom_real_data[224] = -91;
            rom_real_data[225] = -97;
            rom_real_data[226] = -103;
            rom_real_data[227] = -108;
            rom_real_data[228] = -113;
            rom_real_data[229] = -117;
            rom_real_data[230] = -121;
            rom_real_data[231] = -123;
            rom_real_data[232] = -126;
            rom_real_data[233] = -127;
            rom_real_data[234] = -128;
            rom_real_data[235] = -128;
            rom_real_data[236] = -127;
            rom_real_data[237] = -126;
            rom_real_data[238] = -124;
            rom_real_data[239] = -122;
            rom_real_data[240] = -118;
            rom_real_data[241] = -114;
            rom_real_data[242] = -110;
            rom_real_data[243] = -105;
            rom_real_data[244] = -99;
            rom_real_data[245] = -93;
            rom_real_data[246] = -86;
            rom_real_data[247] = -79;
            rom_real_data[248] = -71;
            rom_real_data[249] = -63;
            rom_real_data[250] = -55;
            rom_real_data[251] = -46;
            rom_real_data[252] = -37;
            rom_real_data[253] = -28;
            rom_real_data[254] = -19;
            rom_real_data[255] = -9;
            rom_real_data[256] = 128;
            rom_real_data[257] = 128;
            rom_real_data[258] = 128;
            rom_real_data[259] = 128;
            rom_real_data[260] = 128;
            rom_real_data[261] = 128;
            rom_real_data[262] = 128;
            rom_real_data[263] = 128;
            rom_real_data[264] = 127;
            rom_real_data[265] = 127;
            rom_real_data[266] = 127;
            rom_real_data[267] = 127;
            rom_real_data[268] = 127;
            rom_real_data[269] = 126;
            rom_real_data[270] = 126;
            rom_real_data[271] = 126;
            rom_real_data[272] = 126;
            rom_real_data[273] = 125;
            rom_real_data[274] = 125;
            rom_real_data[275] = 125;
            rom_real_data[276] = 124;
            rom_real_data[277] = 124;
            rom_real_data[278] = 123;
            rom_real_data[279] = 123;
            rom_real_data[280] = 122;
            rom_real_data[281] = 122;
            rom_real_data[282] = 122;
            rom_real_data[283] = 121;
            rom_real_data[284] = 121;
            rom_real_data[285] = 120;
            rom_real_data[286] = 119;
            rom_real_data[287] = 119;
            rom_real_data[288] = 118;
            rom_real_data[289] = 118;
            rom_real_data[290] = 117;
            rom_real_data[291] = 116;
            rom_real_data[292] = 116;
            rom_real_data[293] = 115;
            rom_real_data[294] = 114;
            rom_real_data[295] = 114;
            rom_real_data[296] = 113;
            rom_real_data[297] = 112;
            rom_real_data[298] = 111;
            rom_real_data[299] = 111;
            rom_real_data[300] = 110;
            rom_real_data[301] = 109;
            rom_real_data[302] = 108;
            rom_real_data[303] = 107;
            rom_real_data[304] = 106;
            rom_real_data[305] = 106;
            rom_real_data[306] = 105;
            rom_real_data[307] = 104;
            rom_real_data[308] = 103;
            rom_real_data[309] = 102;
            rom_real_data[310] = 101;
            rom_real_data[311] = 100;
            rom_real_data[312] = 99;
            rom_real_data[313] = 98;
            rom_real_data[314] = 97;
            rom_real_data[315] = 96;
            rom_real_data[316] = 95;
            rom_real_data[317] = 94;
            rom_real_data[318] = 93;
            rom_real_data[319] = 92;
            rom_real_data[320] = 128;
            rom_real_data[321] = 128;
            rom_real_data[322] = 127;
            rom_real_data[323] = 126;
            rom_real_data[324] = 124;
            rom_real_data[325] = 122;
            rom_real_data[326] = 119;
            rom_real_data[327] = 116;
            rom_real_data[328] = 113;
            rom_real_data[329] = 109;
            rom_real_data[330] = 105;
            rom_real_data[331] = 100;
            rom_real_data[332] = 95;
            rom_real_data[333] = 89;
            rom_real_data[334] = 84;
            rom_real_data[335] = 78;
            rom_real_data[336] = 71;
            rom_real_data[337] = 64;
            rom_real_data[338] = 58;
            rom_real_data[339] = 50;
            rom_real_data[340] = 43;
            rom_real_data[341] = 36;
            rom_real_data[342] = 28;
            rom_real_data[343] = 20;
            rom_real_data[344] = 13;
            rom_real_data[345] = 5;
            rom_real_data[346] = -3;
            rom_real_data[347] = -11;
            rom_real_data[348] = -19;
            rom_real_data[349] = -27;
            rom_real_data[350] = -34;
            rom_real_data[351] = -42;
            rom_real_data[352] = -49;
            rom_real_data[353] = -56;
            rom_real_data[354] = -63;
            rom_real_data[355] = -70;
            rom_real_data[356] = -76;
            rom_real_data[357] = -82;
            rom_real_data[358] = -88;
            rom_real_data[359] = -94;
            rom_real_data[360] = -99;
            rom_real_data[361] = -104;
            rom_real_data[362] = -108;
            rom_real_data[363] = -112;
            rom_real_data[364] = -116;
            rom_real_data[365] = -119;
            rom_real_data[366] = -122;
            rom_real_data[367] = -124;
            rom_real_data[368] = -126;
            rom_real_data[369] = -127;
            rom_real_data[370] = -128;
            rom_real_data[371] = -128;
            rom_real_data[372] = -128;
            rom_real_data[373] = -127;
            rom_real_data[374] = -126;
            rom_real_data[375] = -125;
            rom_real_data[376] = -122;
            rom_real_data[377] = -120;
            rom_real_data[378] = -117;
            rom_real_data[379] = -114;
            rom_real_data[380] = -110;
            rom_real_data[381] = -106;
            rom_real_data[382] = -101;
            rom_real_data[383] = -96;
            rom_real_data[384] = 128;
            rom_real_data[385] = 128;
            rom_real_data[386] = 128;
            rom_real_data[387] = 127;
            rom_real_data[388] = 127;
            rom_real_data[389] = 126;
            rom_real_data[390] = 125;
            rom_real_data[391] = 124;
            rom_real_data[392] = 122;
            rom_real_data[393] = 121;
            rom_real_data[394] = 119;
            rom_real_data[395] = 118;
            rom_real_data[396] = 116;
            rom_real_data[397] = 114;
            rom_real_data[398] = 111;
            rom_real_data[399] = 109;
            rom_real_data[400] = 106;
            rom_real_data[401] = 104;
            rom_real_data[402] = 101;
            rom_real_data[403] = 98;
            rom_real_data[404] = 95;
            rom_real_data[405] = 92;
            rom_real_data[406] = 88;
            rom_real_data[407] = 85;
            rom_real_data[408] = 81;
            rom_real_data[409] = 78;
            rom_real_data[410] = 74;
            rom_real_data[411] = 70;
            rom_real_data[412] = 66;
            rom_real_data[413] = 62;
            rom_real_data[414] = 58;
            rom_real_data[415] = 53;
            rom_real_data[416] = 49;
            rom_real_data[417] = 45;
            rom_real_data[418] = 40;
            rom_real_data[419] = 36;
            rom_real_data[420] = 31;
            rom_real_data[421] = 27;
            rom_real_data[422] = 22;
            rom_real_data[423] = 17;
            rom_real_data[424] = 13;
            rom_real_data[425] = 8;
            rom_real_data[426] = 3;
            rom_real_data[427] = -2;
            rom_real_data[428] = -6;
            rom_real_data[429] = -11;
            rom_real_data[430] = -16;
            rom_real_data[431] = -20;
            rom_real_data[432] = -25;
            rom_real_data[433] = -30;
            rom_real_data[434] = -34;
            rom_real_data[435] = -39;
            rom_real_data[436] = -43;
            rom_real_data[437] = -48;
            rom_real_data[438] = -52;
            rom_real_data[439] = -56;
            rom_real_data[440] = -60;
            rom_real_data[441] = -64;
            rom_real_data[442] = -68;
            rom_real_data[443] = -72;
            rom_real_data[444] = -76;
            rom_real_data[445] = -80;
            rom_real_data[446] = -84;
            rom_real_data[447] = -87;
            rom_real_data[448] = 128;
            rom_real_data[449] = 128;
            rom_real_data[450] = 126;
            rom_real_data[451] = 124;
            rom_real_data[452] = 121;
            rom_real_data[453] = 116;
            rom_real_data[454] = 111;
            rom_real_data[455] = 106;
            rom_real_data[456] = 99;
            rom_real_data[457] = 92;
            rom_real_data[458] = 84;
            rom_real_data[459] = 75;
            rom_real_data[460] = 66;
            rom_real_data[461] = 56;
            rom_real_data[462] = 46;
            rom_real_data[463] = 36;
            rom_real_data[464] = 25;
            rom_real_data[465] = 14;
            rom_real_data[466] = 3;
            rom_real_data[467] = -8;
            rom_real_data[468] = -19;
            rom_real_data[469] = -30;
            rom_real_data[470] = -40;
            rom_real_data[471] = -50;
            rom_real_data[472] = -60;
            rom_real_data[473] = -70;
            rom_real_data[474] = -79;
            rom_real_data[475] = -87;
            rom_real_data[476] = -95;
            rom_real_data[477] = -102;
            rom_real_data[478] = -108;
            rom_real_data[479] = -114;
            rom_real_data[480] = -118;
            rom_real_data[481] = -122;
            rom_real_data[482] = -125;
            rom_real_data[483] = -127;
            rom_real_data[484] = -128;
            rom_real_data[485] = -128;
            rom_real_data[486] = -127;
            rom_real_data[487] = -125;
            rom_real_data[488] = -122;
            rom_real_data[489] = -119;
            rom_real_data[490] = -114;
            rom_real_data[491] = -109;
            rom_real_data[492] = -103;
            rom_real_data[493] = -96;
            rom_real_data[494] = -88;
            rom_real_data[495] = -80;
            rom_real_data[496] = -71;
            rom_real_data[497] = -62;
            rom_real_data[498] = -52;
            rom_real_data[499] = -42;
            rom_real_data[500] = -31;
            rom_real_data[501] = -20;
            rom_real_data[502] = -9;
            rom_real_data[503] = 2;
            rom_real_data[504] = 13;
            rom_real_data[505] = 23;
            rom_real_data[506] = 34;
            rom_real_data[507] = 45;
            rom_real_data[508] = 55;
            rom_real_data[509] = 64;
            rom_real_data[510] = 74;
            rom_real_data[511] = 82;




            rom_imag_data[0] = 0;
            rom_imag_data[1] = 0;
            rom_imag_data[2] = 0;
            rom_imag_data[3] = 0;
            rom_imag_data[4] = 0;
            rom_imag_data[5] = 0;
            rom_imag_data[6] = 0;
            rom_imag_data[7] = 0;
            rom_imag_data[8] = 0;
            rom_imag_data[9] = 0;
            rom_imag_data[10] = 0;
            rom_imag_data[11] = 0;
            rom_imag_data[12] = 0;
            rom_imag_data[13] = 0;
            rom_imag_data[14] = 0;
            rom_imag_data[15] = 0;
            rom_imag_data[16] = 0;
            rom_imag_data[17] = 0;
            rom_imag_data[18] = 0;
            rom_imag_data[19] = 0;
            rom_imag_data[20] = 0;
            rom_imag_data[21] = 0;
            rom_imag_data[22] = 0;
            rom_imag_data[23] = 0;
            rom_imag_data[24] = 0;
            rom_imag_data[25] = 0;
            rom_imag_data[26] = 0;
            rom_imag_data[27] = 0;
            rom_imag_data[28] = 0;
            rom_imag_data[29] = 0;
            rom_imag_data[30] = 0;
            rom_imag_data[31] = 0;
            rom_imag_data[32] = 0;
            rom_imag_data[33] = 0;
            rom_imag_data[34] = 0;
            rom_imag_data[35] = 0;
            rom_imag_data[36] = 0;
            rom_imag_data[37] = 0;
            rom_imag_data[38] = 0;
            rom_imag_data[39] = 0;
            rom_imag_data[40] = 0;
            rom_imag_data[41] = 0;
            rom_imag_data[42] = 0;
            rom_imag_data[43] = 0;
            rom_imag_data[44] = 0;
            rom_imag_data[45] = 0;
            rom_imag_data[46] = 0;
            rom_imag_data[47] = 0;
            rom_imag_data[48] = 0;
            rom_imag_data[49] = 0;
            rom_imag_data[50] = 0;
            rom_imag_data[51] = 0;
            rom_imag_data[52] = 0;
            rom_imag_data[53] = 0;
            rom_imag_data[54] = 0;
            rom_imag_data[55] = 0;
            rom_imag_data[56] = 0;
            rom_imag_data[57] = 0;
            rom_imag_data[58] = 0;
            rom_imag_data[59] = 0;
            rom_imag_data[60] = 0;
            rom_imag_data[61] = 0;
            rom_imag_data[62] = 0;
            rom_imag_data[63] = 0;
            rom_imag_data[64] = 0;
            rom_imag_data[65] = -6;
            rom_imag_data[66] = -13;
            rom_imag_data[67] = -19;
            rom_imag_data[68] = -25;
            rom_imag_data[69] = -31;
            rom_imag_data[70] = -37;
            rom_imag_data[71] = -43;
            rom_imag_data[72] = -49;
            rom_imag_data[73] = -55;
            rom_imag_data[74] = -60;
            rom_imag_data[75] = -66;
            rom_imag_data[76] = -71;
            rom_imag_data[77] = -76;
            rom_imag_data[78] = -81;
            rom_imag_data[79] = -86;
            rom_imag_data[80] = -91;
            rom_imag_data[81] = -95;
            rom_imag_data[82] = -99;
            rom_imag_data[83] = -103;
            rom_imag_data[84] = -106;
            rom_imag_data[85] = -110;
            rom_imag_data[86] = -113;
            rom_imag_data[87] = -116;
            rom_imag_data[88] = -118;
            rom_imag_data[89] = -121;
            rom_imag_data[90] = -122;
            rom_imag_data[91] = -124;
            rom_imag_data[92] = -126;
            rom_imag_data[93] = -127;
            rom_imag_data[94] = -127;
            rom_imag_data[95] = -128;
            rom_imag_data[96] = -128;
            rom_imag_data[97] = -128;
            rom_imag_data[98] = -127;
            rom_imag_data[99] = -127;
            rom_imag_data[100] = -126;
            rom_imag_data[101] = -124;
            rom_imag_data[102] = -122;
            rom_imag_data[103] = -121;
            rom_imag_data[104] = -118;
            rom_imag_data[105] = -116;
            rom_imag_data[106] = -113;
            rom_imag_data[107] = -110;
            rom_imag_data[108] = -106;
            rom_imag_data[109] = -103;
            rom_imag_data[110] = -99;
            rom_imag_data[111] = -95;
            rom_imag_data[112] = -91;
            rom_imag_data[113] = -86;
            rom_imag_data[114] = -81;
            rom_imag_data[115] = -76;
            rom_imag_data[116] = -71;
            rom_imag_data[117] = -66;
            rom_imag_data[118] = -60;
            rom_imag_data[119] = -55;
            rom_imag_data[120] = -49;
            rom_imag_data[121] = -43;
            rom_imag_data[122] = -37;
            rom_imag_data[123] = -31;
            rom_imag_data[124] = -25;
            rom_imag_data[125] = -19;
            rom_imag_data[126] = -13;
            rom_imag_data[127] = -6;
            rom_imag_data[128] = 0;
            rom_imag_data[129] = -3;
            rom_imag_data[130] = -6;
            rom_imag_data[131] = -9;
            rom_imag_data[132] = -13;
            rom_imag_data[133] = -16;
            rom_imag_data[134] = -19;
            rom_imag_data[135] = -22;
            rom_imag_data[136] = -25;
            rom_imag_data[137] = -28;
            rom_imag_data[138] = -31;
            rom_imag_data[139] = -34;
            rom_imag_data[140] = -37;
            rom_imag_data[141] = -40;
            rom_imag_data[142] = -43;
            rom_imag_data[143] = -46;
            rom_imag_data[144] = -49;
            rom_imag_data[145] = -52;
            rom_imag_data[146] = -55;
            rom_imag_data[147] = -58;
            rom_imag_data[148] = -60;
            rom_imag_data[149] = -63;
            rom_imag_data[150] = -66;
            rom_imag_data[151] = -68;
            rom_imag_data[152] = -71;
            rom_imag_data[153] = -74;
            rom_imag_data[154] = -76;
            rom_imag_data[155] = -79;
            rom_imag_data[156] = -81;
            rom_imag_data[157] = -84;
            rom_imag_data[158] = -86;
            rom_imag_data[159] = -88;
            rom_imag_data[160] = -91;
            rom_imag_data[161] = -93;
            rom_imag_data[162] = -95;
            rom_imag_data[163] = -97;
            rom_imag_data[164] = -99;
            rom_imag_data[165] = -101;
            rom_imag_data[166] = -103;
            rom_imag_data[167] = -105;
            rom_imag_data[168] = -106;
            rom_imag_data[169] = -108;
            rom_imag_data[170] = -110;
            rom_imag_data[171] = -111;
            rom_imag_data[172] = -113;
            rom_imag_data[173] = -114;
            rom_imag_data[174] = -116;
            rom_imag_data[175] = -117;
            rom_imag_data[176] = -118;
            rom_imag_data[177] = -119;
            rom_imag_data[178] = -121;
            rom_imag_data[179] = -122;
            rom_imag_data[180] = -122;
            rom_imag_data[181] = -123;
            rom_imag_data[182] = -124;
            rom_imag_data[183] = -125;
            rom_imag_data[184] = -126;
            rom_imag_data[185] = -126;
            rom_imag_data[186] = -127;
            rom_imag_data[187] = -127;
            rom_imag_data[188] = -127;
            rom_imag_data[189] = -128;
            rom_imag_data[190] = -128;
            rom_imag_data[191] = -128;
            rom_imag_data[192] = 0;
            rom_imag_data[193] = -9;
            rom_imag_data[194] = -19;
            rom_imag_data[195] = -28;
            rom_imag_data[196] = -37;
            rom_imag_data[197] = -46;
            rom_imag_data[198] = -55;
            rom_imag_data[199] = -63;
            rom_imag_data[200] = -71;
            rom_imag_data[201] = -79;
            rom_imag_data[202] = -86;
            rom_imag_data[203] = -93;
            rom_imag_data[204] = -99;
            rom_imag_data[205] = -105;
            rom_imag_data[206] = -110;
            rom_imag_data[207] = -114;
            rom_imag_data[208] = -118;
            rom_imag_data[209] = -122;
            rom_imag_data[210] = -124;
            rom_imag_data[211] = -126;
            rom_imag_data[212] = -127;
            rom_imag_data[213] = -128;
            rom_imag_data[214] = -128;
            rom_imag_data[215] = -127;
            rom_imag_data[216] = -126;
            rom_imag_data[217] = -123;
            rom_imag_data[218] = -121;
            rom_imag_data[219] = -117;
            rom_imag_data[220] = -113;
            rom_imag_data[221] = -108;
            rom_imag_data[222] = -103;
            rom_imag_data[223] = -97;
            rom_imag_data[224] = -91;
            rom_imag_data[225] = -84;
            rom_imag_data[226] = -76;
            rom_imag_data[227] = -68;
            rom_imag_data[228] = -60;
            rom_imag_data[229] = -52;
            rom_imag_data[230] = -43;
            rom_imag_data[231] = -34;
            rom_imag_data[232] = -25;
            rom_imag_data[233] = -16;
            rom_imag_data[234] = -6;
            rom_imag_data[235] = 3;
            rom_imag_data[236] = 13;
            rom_imag_data[237] = 22;
            rom_imag_data[238] = 31;
            rom_imag_data[239] = 40;
            rom_imag_data[240] = 49;
            rom_imag_data[241] = 58;
            rom_imag_data[242] = 66;
            rom_imag_data[243] = 74;
            rom_imag_data[244] = 81;
            rom_imag_data[245] = 88;
            rom_imag_data[246] = 95;
            rom_imag_data[247] = 101;
            rom_imag_data[248] = 106;
            rom_imag_data[249] = 111;
            rom_imag_data[250] = 116;
            rom_imag_data[251] = 119;
            rom_imag_data[252] = 122;
            rom_imag_data[253] = 125;
            rom_imag_data[254] = 127;
            rom_imag_data[255] = 128;
            rom_imag_data[256] = 0;
            rom_imag_data[257] = -2;
            rom_imag_data[258] = -3;
            rom_imag_data[259] = -5;
            rom_imag_data[260] = -6;
            rom_imag_data[261] = -8;
            rom_imag_data[262] = -9;
            rom_imag_data[263] = -11;
            rom_imag_data[264] = -13;
            rom_imag_data[265] = -14;
            rom_imag_data[266] = -16;
            rom_imag_data[267] = -17;
            rom_imag_data[268] = -19;
            rom_imag_data[269] = -20;
            rom_imag_data[270] = -22;
            rom_imag_data[271] = -23;
            rom_imag_data[272] = -25;
            rom_imag_data[273] = -27;
            rom_imag_data[274] = -28;
            rom_imag_data[275] = -30;
            rom_imag_data[276] = -31;
            rom_imag_data[277] = -33;
            rom_imag_data[278] = -34;
            rom_imag_data[279] = -36;
            rom_imag_data[280] = -37;
            rom_imag_data[281] = -39;
            rom_imag_data[282] = -40;
            rom_imag_data[283] = -42;
            rom_imag_data[284] = -43;
            rom_imag_data[285] = -45;
            rom_imag_data[286] = -46;
            rom_imag_data[287] = -48;
            rom_imag_data[288] = -49;
            rom_imag_data[289] = -50;
            rom_imag_data[290] = -52;
            rom_imag_data[291] = -53;
            rom_imag_data[292] = -55;
            rom_imag_data[293] = -56;
            rom_imag_data[294] = -58;
            rom_imag_data[295] = -59;
            rom_imag_data[296] = -60;
            rom_imag_data[297] = -62;
            rom_imag_data[298] = -63;
            rom_imag_data[299] = -64;
            rom_imag_data[300] = -66;
            rom_imag_data[301] = -67;
            rom_imag_data[302] = -68;
            rom_imag_data[303] = -70;
            rom_imag_data[304] = -71;
            rom_imag_data[305] = -72;
            rom_imag_data[306] = -74;
            rom_imag_data[307] = -75;
            rom_imag_data[308] = -76;
            rom_imag_data[309] = -78;
            rom_imag_data[310] = -79;
            rom_imag_data[311] = -80;
            rom_imag_data[312] = -81;
            rom_imag_data[313] = -82;
            rom_imag_data[314] = -84;
            rom_imag_data[315] = -85;
            rom_imag_data[316] = -86;
            rom_imag_data[317] = -87;
            rom_imag_data[318] = -88;
            rom_imag_data[319] = -89;
            rom_imag_data[320] = 0;
            rom_imag_data[321] = -8;
            rom_imag_data[322] = -16;
            rom_imag_data[323] = -23;
            rom_imag_data[324] = -31;
            rom_imag_data[325] = -39;
            rom_imag_data[326] = -46;
            rom_imag_data[327] = -53;
            rom_imag_data[328] = -60;
            rom_imag_data[329] = -67;
            rom_imag_data[330] = -74;
            rom_imag_data[331] = -80;
            rom_imag_data[332] = -86;
            rom_imag_data[333] = -92;
            rom_imag_data[334] = -97;
            rom_imag_data[335] = -102;
            rom_imag_data[336] = -106;
            rom_imag_data[337] = -111;
            rom_imag_data[338] = -114;
            rom_imag_data[339] = -118;
            rom_imag_data[340] = -121;
            rom_imag_data[341] = -123;
            rom_imag_data[342] = -125;
            rom_imag_data[343] = -126;
            rom_imag_data[344] = -127;
            rom_imag_data[345] = -128;
            rom_imag_data[346] = -128;
            rom_imag_data[347] = -128;
            rom_imag_data[348] = -127;
            rom_imag_data[349] = -125;
            rom_imag_data[350] = -123;
            rom_imag_data[351] = -121;
            rom_imag_data[352] = -118;
            rom_imag_data[353] = -115;
            rom_imag_data[354] = -111;
            rom_imag_data[355] = -107;
            rom_imag_data[356] = -103;
            rom_imag_data[357] = -98;
            rom_imag_data[358] = -93;
            rom_imag_data[359] = -87;
            rom_imag_data[360] = -81;
            rom_imag_data[361] = -75;
            rom_imag_data[362] = -68;
            rom_imag_data[363] = -62;
            rom_imag_data[364] = -55;
            rom_imag_data[365] = -48;
            rom_imag_data[366] = -40;
            rom_imag_data[367] = -33;
            rom_imag_data[368] = -25;
            rom_imag_data[369] = -17;
            rom_imag_data[370] = -9;
            rom_imag_data[371] = -2;
            rom_imag_data[372] = 6;
            rom_imag_data[373] = 14;
            rom_imag_data[374] = 22;
            rom_imag_data[375] = 30;
            rom_imag_data[376] = 37;
            rom_imag_data[377] = 45;
            rom_imag_data[378] = 52;
            rom_imag_data[379] = 59;
            rom_imag_data[380] = 66;
            rom_imag_data[381] = 72;
            rom_imag_data[382] = 79;
            rom_imag_data[383] = 85;
            rom_imag_data[384] = 0;
            rom_imag_data[385] = -5;
            rom_imag_data[386] = -9;
            rom_imag_data[387] = -14;
            rom_imag_data[388] = -19;
            rom_imag_data[389] = -23;
            rom_imag_data[390] = -28;
            rom_imag_data[391] = -33;
            rom_imag_data[392] = -37;
            rom_imag_data[393] = -42;
            rom_imag_data[394] = -46;
            rom_imag_data[395] = -50;
            rom_imag_data[396] = -55;
            rom_imag_data[397] = -59;
            rom_imag_data[398] = -63;
            rom_imag_data[399] = -67;
            rom_imag_data[400] = -71;
            rom_imag_data[401] = -75;
            rom_imag_data[402] = -79;
            rom_imag_data[403] = -82;
            rom_imag_data[404] = -86;
            rom_imag_data[405] = -89;
            rom_imag_data[406] = -93;
            rom_imag_data[407] = -96;
            rom_imag_data[408] = -99;
            rom_imag_data[409] = -102;
            rom_imag_data[410] = -105;
            rom_imag_data[411] = -107;
            rom_imag_data[412] = -110;
            rom_imag_data[413] = -112;
            rom_imag_data[414] = -114;
            rom_imag_data[415] = -116;
            rom_imag_data[416] = -118;
            rom_imag_data[417] = -120;
            rom_imag_data[418] = -122;
            rom_imag_data[419] = -123;
            rom_imag_data[420] = -124;
            rom_imag_data[421] = -125;
            rom_imag_data[422] = -126;
            rom_imag_data[423] = -127;
            rom_imag_data[424] = -127;
            rom_imag_data[425] = -128;
            rom_imag_data[426] = -128;
            rom_imag_data[427] = -128;
            rom_imag_data[428] = -128;
            rom_imag_data[429] = -128;
            rom_imag_data[430] = -127;
            rom_imag_data[431] = -126;
            rom_imag_data[432] = -126;
            rom_imag_data[433] = -125;
            rom_imag_data[434] = -123;
            rom_imag_data[435] = -122;
            rom_imag_data[436] = -121;
            rom_imag_data[437] = -119;
            rom_imag_data[438] = -117;
            rom_imag_data[439] = -115;
            rom_imag_data[440] = -113;
            rom_imag_data[441] = -111;
            rom_imag_data[442] = -108;
            rom_imag_data[443] = -106;
            rom_imag_data[444] = -103;
            rom_imag_data[445] = -100;
            rom_imag_data[446] = -97;
            rom_imag_data[447] = -94;
            rom_imag_data[448] = 0;
            rom_imag_data[449] = -11;
            rom_imag_data[450] = -22;
            rom_imag_data[451] = -33;
            rom_imag_data[452] = -43;
            rom_imag_data[453] = -53;
            rom_imag_data[454] = -63;
            rom_imag_data[455] = -72;
            rom_imag_data[456] = -81;
            rom_imag_data[457] = -89;
            rom_imag_data[458] = -97;
            rom_imag_data[459] = -104;
            rom_imag_data[460] = -110;
            rom_imag_data[461] = -115;
            rom_imag_data[462] = -119;
            rom_imag_data[463] = -123;
            rom_imag_data[464] = -126;
            rom_imag_data[465] = -127;
            rom_imag_data[466] = -128;
            rom_imag_data[467] = -128;
            rom_imag_data[468] = -127;
            rom_imag_data[469] = -125;
            rom_imag_data[470] = -122;
            rom_imag_data[471] = -118;
            rom_imag_data[472] = -113;
            rom_imag_data[473] = -107;
            rom_imag_data[474] = -101;
            rom_imag_data[475] = -94;
            rom_imag_data[476] = -86;
            rom_imag_data[477] = -78;
            rom_imag_data[478] = -68;
            rom_imag_data[479] = -59;
            rom_imag_data[480] = -49;
            rom_imag_data[481] = -39;
            rom_imag_data[482] = -28;
            rom_imag_data[483] = -17;
            rom_imag_data[484] = -6;
            rom_imag_data[485] = 5;
            rom_imag_data[486] = 16;
            rom_imag_data[487] = 27;
            rom_imag_data[488] = 37;
            rom_imag_data[489] = 48;
            rom_imag_data[490] = 58;
            rom_imag_data[491] = 67;
            rom_imag_data[492] = 76;
            rom_imag_data[493] = 85;
            rom_imag_data[494] = 93;
            rom_imag_data[495] = 100;
            rom_imag_data[496] = 106;
            rom_imag_data[497] = 112;
            rom_imag_data[498] = 117;
            rom_imag_data[499] = 121;
            rom_imag_data[500] = 124;
            rom_imag_data[501] = 126;
            rom_imag_data[502] = 128;
            rom_imag_data[503] = 128;
            rom_imag_data[504] = 127;
            rom_imag_data[505] = 126;
            rom_imag_data[506] = 123;
            rom_imag_data[507] = 120;
            rom_imag_data[508] = 116;
            rom_imag_data[509] = 111;
            rom_imag_data[510] = 105;
            rom_imag_data[511] = 98;
            end
            else begin
                rom_real_data[0] = 128;
            rom_real_data[1] = 128;
            rom_real_data[2] = 128;
            rom_real_data[3] = 128;
            rom_real_data[4] = 128;
            rom_real_data[5] = 128;
            rom_real_data[6] = 128;
            rom_real_data[7] = 128;
            rom_real_data[8] = 128;
            rom_real_data[9] = 128;
            rom_real_data[10] = 128;
            rom_real_data[11] = 128;
            rom_real_data[12] = 128;
            rom_real_data[13] = 128;
            rom_real_data[14] = 128;
            rom_real_data[15] = 128;
            rom_real_data[16] = 128;
            rom_real_data[17] = 128;
            rom_real_data[18] = 128;
            rom_real_data[19] = 128;
            rom_real_data[20] = 128;
            rom_real_data[21] = 128;
            rom_real_data[22] = 128;
            rom_real_data[23] = 128;
            rom_real_data[24] = 128;
            rom_real_data[25] = 128;
            rom_real_data[26] = 128;
            rom_real_data[27] = 128;
            rom_real_data[28] = 128;
            rom_real_data[29] = 128;
            rom_real_data[30] = 128;
            rom_real_data[31] = 128;
            rom_real_data[32] = 128;
            rom_real_data[33] = 128;
            rom_real_data[34] = 128;
            rom_real_data[35] = 128;
            rom_real_data[36] = 128;
            rom_real_data[37] = 128;
            rom_real_data[38] = 128;
            rom_real_data[39] = 128;
            rom_real_data[40] = 128;
            rom_real_data[41] = 128;
            rom_real_data[42] = 128;
            rom_real_data[43] = 128;
            rom_real_data[44] = 128;
            rom_real_data[45] = 128;
            rom_real_data[46] = 128;
            rom_real_data[47] = 128;
            rom_real_data[48] = 128;
            rom_real_data[49] = 128;
            rom_real_data[50] = 128;
            rom_real_data[51] = 128;
            rom_real_data[52] = 128;
            rom_real_data[53] = 128;
            rom_real_data[54] = 128;
            rom_real_data[55] = 128;
            rom_real_data[56] = 128;
            rom_real_data[57] = 128;
            rom_real_data[58] = 128;
            rom_real_data[59] = 128;
            rom_real_data[60] = 128;
            rom_real_data[61] = 128;
            rom_real_data[62] = 128;
            rom_real_data[63] = 128;
            rom_real_data[64] = 128;
            rom_real_data[65] = 128;
            rom_real_data[66] = 127;
            rom_real_data[67] = 127;
            rom_real_data[68] = 126;
            rom_real_data[69] = 124;
            rom_real_data[70] = 122;
            rom_real_data[71] = 121;
            rom_real_data[72] = 118;
            rom_real_data[73] = 116;
            rom_real_data[74] = 113;
            rom_real_data[75] = 110;
            rom_real_data[76] = 106;
            rom_real_data[77] = 103;
            rom_real_data[78] = 99;
            rom_real_data[79] = 95;
            rom_real_data[80] = 91;
            rom_real_data[81] = 86;
            rom_real_data[82] = 81;
            rom_real_data[83] = 76;
            rom_real_data[84] = 71;
            rom_real_data[85] = 66;
            rom_real_data[86] = 60;
            rom_real_data[87] = 55;
            rom_real_data[88] = 49;
            rom_real_data[89] = 43;
            rom_real_data[90] = 37;
            rom_real_data[91] = 31;
            rom_real_data[92] = 25;
            rom_real_data[93] = 19;
            rom_real_data[94] = 13;
            rom_real_data[95] = 6;
            rom_real_data[96] = 0;
            rom_real_data[97] = -6;
            rom_real_data[98] = -13;
            rom_real_data[99] = -19;
            rom_real_data[100] = -25;
            rom_real_data[101] = -31;
            rom_real_data[102] = -37;
            rom_real_data[103] = -43;
            rom_real_data[104] = -49;
            rom_real_data[105] = -55;
            rom_real_data[106] = -60;
            rom_real_data[107] = -66;
            rom_real_data[108] = -71;
            rom_real_data[109] = -76;
            rom_real_data[110] = -81;
            rom_real_data[111] = -86;
            rom_real_data[112] = -91;
            rom_real_data[113] = -95;
            rom_real_data[114] = -99;
            rom_real_data[115] = -103;
            rom_real_data[116] = -106;
            rom_real_data[117] = -110;
            rom_real_data[118] = -113;
            rom_real_data[119] = -116;
            rom_real_data[120] = -118;
            rom_real_data[121] = -121;
            rom_real_data[122] = -122;
            rom_real_data[123] = -124;
            rom_real_data[124] = -126;
            rom_real_data[125] = -127;
            rom_real_data[126] = -127;
            rom_real_data[127] = -128;
            rom_real_data[128] = 128;
            rom_real_data[129] = 128;
            rom_real_data[130] = 128;
            rom_real_data[131] = 128;
            rom_real_data[132] = 127;
            rom_real_data[133] = 127;
            rom_real_data[134] = 127;
            rom_real_data[135] = 126;
            rom_real_data[136] = 126;
            rom_real_data[137] = 125;
            rom_real_data[138] = 124;
            rom_real_data[139] = 123;
            rom_real_data[140] = 122;
            rom_real_data[141] = 122;
            rom_real_data[142] = 121;
            rom_real_data[143] = 119;
            rom_real_data[144] = 118;
            rom_real_data[145] = 117;
            rom_real_data[146] = 116;
            rom_real_data[147] = 114;
            rom_real_data[148] = 113;
            rom_real_data[149] = 111;
            rom_real_data[150] = 110;
            rom_real_data[151] = 108;
            rom_real_data[152] = 106;
            rom_real_data[153] = 105;
            rom_real_data[154] = 103;
            rom_real_data[155] = 101;
            rom_real_data[156] = 99;
            rom_real_data[157] = 97;
            rom_real_data[158] = 95;
            rom_real_data[159] = 93;
            rom_real_data[160] = 91;
            rom_real_data[161] = 88;
            rom_real_data[162] = 86;
            rom_real_data[163] = 84;
            rom_real_data[164] = 81;
            rom_real_data[165] = 79;
            rom_real_data[166] = 76;
            rom_real_data[167] = 74;
            rom_real_data[168] = 71;
            rom_real_data[169] = 68;
            rom_real_data[170] = 66;
            rom_real_data[171] = 63;
            rom_real_data[172] = 60;
            rom_real_data[173] = 58;
            rom_real_data[174] = 55;
            rom_real_data[175] = 52;
            rom_real_data[176] = 49;
            rom_real_data[177] = 46;
            rom_real_data[178] = 43;
            rom_real_data[179] = 40;
            rom_real_data[180] = 37;
            rom_real_data[181] = 34;
            rom_real_data[182] = 31;
            rom_real_data[183] = 28;
            rom_real_data[184] = 25;
            rom_real_data[185] = 22;
            rom_real_data[186] = 19;
            rom_real_data[187] = 16;
            rom_real_data[188] = 13;
            rom_real_data[189] = 9;
            rom_real_data[190] = 6;
            rom_real_data[191] = 3;
            rom_real_data[192] = 128;
            rom_real_data[193] = 128;
            rom_real_data[194] = 127;
            rom_real_data[195] = 125;
            rom_real_data[196] = 122;
            rom_real_data[197] = 119;
            rom_real_data[198] = 116;
            rom_real_data[199] = 111;
            rom_real_data[200] = 106;
            rom_real_data[201] = 101;
            rom_real_data[202] = 95;
            rom_real_data[203] = 88;
            rom_real_data[204] = 81;
            rom_real_data[205] = 74;
            rom_real_data[206] = 66;
            rom_real_data[207] = 58;
            rom_real_data[208] = 49;
            rom_real_data[209] = 40;
            rom_real_data[210] = 31;
            rom_real_data[211] = 22;
            rom_real_data[212] = 13;
            rom_real_data[213] = 3;
            rom_real_data[214] = -6;
            rom_real_data[215] = -16;
            rom_real_data[216] = -25;
            rom_real_data[217] = -34;
            rom_real_data[218] = -43;
            rom_real_data[219] = -52;
            rom_real_data[220] = -60;
            rom_real_data[221] = -68;
            rom_real_data[222] = -76;
            rom_real_data[223] = -84;
            rom_real_data[224] = -91;
            rom_real_data[225] = -97;
            rom_real_data[226] = -103;
            rom_real_data[227] = -108;
            rom_real_data[228] = -113;
            rom_real_data[229] = -117;
            rom_real_data[230] = -121;
            rom_real_data[231] = -123;
            rom_real_data[232] = -126;
            rom_real_data[233] = -127;
            rom_real_data[234] = -128;
            rom_real_data[235] = -128;
            rom_real_data[236] = -127;
            rom_real_data[237] = -126;
            rom_real_data[238] = -124;
            rom_real_data[239] = -122;
            rom_real_data[240] = -118;
            rom_real_data[241] = -114;
            rom_real_data[242] = -110;
            rom_real_data[243] = -105;
            rom_real_data[244] = -99;
            rom_real_data[245] = -93;
            rom_real_data[246] = -86;
            rom_real_data[247] = -79;
            rom_real_data[248] = -71;
            rom_real_data[249] = -63;
            rom_real_data[250] = -55;
            rom_real_data[251] = -46;
            rom_real_data[252] = -37;
            rom_real_data[253] = -28;
            rom_real_data[254] = -19;
            rom_real_data[255] = -9;
            rom_real_data[256] = 128;
            rom_real_data[257] = 128;
            rom_real_data[258] = 128;
            rom_real_data[259] = 128;
            rom_real_data[260] = 128;
            rom_real_data[261] = 128;
            rom_real_data[262] = 128;
            rom_real_data[263] = 128;
            rom_real_data[264] = 127;
            rom_real_data[265] = 127;
            rom_real_data[266] = 127;
            rom_real_data[267] = 127;
            rom_real_data[268] = 127;
            rom_real_data[269] = 126;
            rom_real_data[270] = 126;
            rom_real_data[271] = 126;
            rom_real_data[272] = 126;
            rom_real_data[273] = 125;
            rom_real_data[274] = 125;
            rom_real_data[275] = 125;
            rom_real_data[276] = 124;
            rom_real_data[277] = 124;
            rom_real_data[278] = 123;
            rom_real_data[279] = 123;
            rom_real_data[280] = 122;
            rom_real_data[281] = 122;
            rom_real_data[282] = 122;
            rom_real_data[283] = 121;
            rom_real_data[284] = 121;
            rom_real_data[285] = 120;
            rom_real_data[286] = 119;
            rom_real_data[287] = 119;
            rom_real_data[288] = 118;
            rom_real_data[289] = 118;
            rom_real_data[290] = 117;
            rom_real_data[291] = 116;
            rom_real_data[292] = 116;
            rom_real_data[293] = 115;
            rom_real_data[294] = 114;
            rom_real_data[295] = 114;
            rom_real_data[296] = 113;
            rom_real_data[297] = 112;
            rom_real_data[298] = 111;
            rom_real_data[299] = 111;
            rom_real_data[300] = 110;
            rom_real_data[301] = 109;
            rom_real_data[302] = 108;
            rom_real_data[303] = 107;
            rom_real_data[304] = 106;
            rom_real_data[305] = 106;
            rom_real_data[306] = 105;
            rom_real_data[307] = 104;
            rom_real_data[308] = 103;
            rom_real_data[309] = 102;
            rom_real_data[310] = 101;
            rom_real_data[311] = 100;
            rom_real_data[312] = 99;
            rom_real_data[313] = 98;
            rom_real_data[314] = 97;
            rom_real_data[315] = 96;
            rom_real_data[316] = 95;
            rom_real_data[317] = 94;
            rom_real_data[318] = 93;
            rom_real_data[319] = 92;
            rom_real_data[320] = 128;
            rom_real_data[321] = 128;
            rom_real_data[322] = 127;
            rom_real_data[323] = 126;
            rom_real_data[324] = 124;
            rom_real_data[325] = 122;
            rom_real_data[326] = 119;
            rom_real_data[327] = 116;
            rom_real_data[328] = 113;
            rom_real_data[329] = 109;
            rom_real_data[330] = 105;
            rom_real_data[331] = 100;
            rom_real_data[332] = 95;
            rom_real_data[333] = 89;
            rom_real_data[334] = 84;
            rom_real_data[335] = 78;
            rom_real_data[336] = 71;
            rom_real_data[337] = 64;
            rom_real_data[338] = 58;
            rom_real_data[339] = 50;
            rom_real_data[340] = 43;
            rom_real_data[341] = 36;
            rom_real_data[342] = 28;
            rom_real_data[343] = 20;
            rom_real_data[344] = 13;
            rom_real_data[345] = 5;
            rom_real_data[346] = -3;
            rom_real_data[347] = -11;
            rom_real_data[348] = -19;
            rom_real_data[349] = -27;
            rom_real_data[350] = -34;
            rom_real_data[351] = -42;
            rom_real_data[352] = -49;
            rom_real_data[353] = -56;
            rom_real_data[354] = -63;
            rom_real_data[355] = -70;
            rom_real_data[356] = -76;
            rom_real_data[357] = -82;
            rom_real_data[358] = -88;
            rom_real_data[359] = -94;
            rom_real_data[360] = -99;
            rom_real_data[361] = -104;
            rom_real_data[362] = -108;
            rom_real_data[363] = -112;
            rom_real_data[364] = -116;
            rom_real_data[365] = -119;
            rom_real_data[366] = -122;
            rom_real_data[367] = -124;
            rom_real_data[368] = -126;
            rom_real_data[369] = -127;
            rom_real_data[370] = -128;
            rom_real_data[371] = -128;
            rom_real_data[372] = -128;
            rom_real_data[373] = -127;
            rom_real_data[374] = -126;
            rom_real_data[375] = -125;
            rom_real_data[376] = -122;
            rom_real_data[377] = -120;
            rom_real_data[378] = -117;
            rom_real_data[379] = -114;
            rom_real_data[380] = -110;
            rom_real_data[381] = -106;
            rom_real_data[382] = -101;
            rom_real_data[383] = -96;
            rom_real_data[384] = 128;
            rom_real_data[385] = 128;
            rom_real_data[386] = 128;
            rom_real_data[387] = 127;
            rom_real_data[388] = 127;
            rom_real_data[389] = 126;
            rom_real_data[390] = 125;
            rom_real_data[391] = 124;
            rom_real_data[392] = 122;
            rom_real_data[393] = 121;
            rom_real_data[394] = 119;
            rom_real_data[395] = 118;
            rom_real_data[396] = 116;
            rom_real_data[397] = 114;
            rom_real_data[398] = 111;
            rom_real_data[399] = 109;
            rom_real_data[400] = 106;
            rom_real_data[401] = 104;
            rom_real_data[402] = 101;
            rom_real_data[403] = 98;
            rom_real_data[404] = 95;
            rom_real_data[405] = 92;
            rom_real_data[406] = 88;
            rom_real_data[407] = 85;
            rom_real_data[408] = 81;
            rom_real_data[409] = 78;
            rom_real_data[410] = 74;
            rom_real_data[411] = 70;
            rom_real_data[412] = 66;
            rom_real_data[413] = 62;
            rom_real_data[414] = 58;
            rom_real_data[415] = 53;
            rom_real_data[416] = 49;
            rom_real_data[417] = 45;
            rom_real_data[418] = 40;
            rom_real_data[419] = 36;
            rom_real_data[420] = 31;
            rom_real_data[421] = 27;
            rom_real_data[422] = 22;
            rom_real_data[423] = 17;
            rom_real_data[424] = 13;
            rom_real_data[425] = 8;
            rom_real_data[426] = 3;
            rom_real_data[427] = -2;
            rom_real_data[428] = -6;
            rom_real_data[429] = -11;
            rom_real_data[430] = -16;
            rom_real_data[431] = -20;
            rom_real_data[432] = -25;
            rom_real_data[433] = -30;
            rom_real_data[434] = -34;
            rom_real_data[435] = -39;
            rom_real_data[436] = -43;
            rom_real_data[437] = -48;
            rom_real_data[438] = -52;
            rom_real_data[439] = -56;
            rom_real_data[440] = -60;
            rom_real_data[441] = -64;
            rom_real_data[442] = -68;
            rom_real_data[443] = -72;
            rom_real_data[444] = -76;
            rom_real_data[445] = -80;
            rom_real_data[446] = -84;
            rom_real_data[447] = -87;
            rom_real_data[448] = 128;
            rom_real_data[449] = 128;
            rom_real_data[450] = 126;
            rom_real_data[451] = 124;
            rom_real_data[452] = 121;
            rom_real_data[453] = 116;
            rom_real_data[454] = 111;
            rom_real_data[455] = 106;
            rom_real_data[456] = 99;
            rom_real_data[457] = 92;
            rom_real_data[458] = 84;
            rom_real_data[459] = 75;
            rom_real_data[460] = 66;
            rom_real_data[461] = 56;
            rom_real_data[462] = 46;
            rom_real_data[463] = 36;
            rom_real_data[464] = 25;
            rom_real_data[465] = 14;
            rom_real_data[466] = 3;
            rom_real_data[467] = -8;
            rom_real_data[468] = -19;
            rom_real_data[469] = -30;
            rom_real_data[470] = -40;
            rom_real_data[471] = -50;
            rom_real_data[472] = -60;
            rom_real_data[473] = -70;
            rom_real_data[474] = -79;
            rom_real_data[475] = -87;
            rom_real_data[476] = -95;
            rom_real_data[477] = -102;
            rom_real_data[478] = -108;
            rom_real_data[479] = -114;
            rom_real_data[480] = -118;
            rom_real_data[481] = -122;
            rom_real_data[482] = -125;
            rom_real_data[483] = -127;
            rom_real_data[484] = -128;
            rom_real_data[485] = -128;
            rom_real_data[486] = -127;
            rom_real_data[487] = -125;
            rom_real_data[488] = -122;
            rom_real_data[489] = -119;
            rom_real_data[490] = -114;
            rom_real_data[491] = -109;
            rom_real_data[492] = -103;
            rom_real_data[493] = -96;
            rom_real_data[494] = -88;
            rom_real_data[495] = -80;
            rom_real_data[496] = -71;
            rom_real_data[497] = -62;
            rom_real_data[498] = -52;
            rom_real_data[499] = -42;
            rom_real_data[500] = -31;
            rom_real_data[501] = -20;
            rom_real_data[502] = -9;
            rom_real_data[503] = 2;
            rom_real_data[504] = 13;
            rom_real_data[505] = 23;
            rom_real_data[506] = 34;
            rom_real_data[507] = 45;
            rom_real_data[508] = 55;
            rom_real_data[509] = 64;
            rom_real_data[510] = 74;
            rom_real_data[511] = 82;




            rom_imag_data[0] = 0;
            rom_imag_data[1] = 0;
            rom_imag_data[2] = 0;
            rom_imag_data[3] = 0;
            rom_imag_data[4] = 0;
            rom_imag_data[5] = 0;
            rom_imag_data[6] = 0;
            rom_imag_data[7] = 0;
            rom_imag_data[8] = 0;
            rom_imag_data[9] = 0;
            rom_imag_data[10] = 0;
            rom_imag_data[11] = 0;
            rom_imag_data[12] = 0;
            rom_imag_data[13] = 0;
            rom_imag_data[14] = 0;
            rom_imag_data[15] = 0;
            rom_imag_data[16] = 0;
            rom_imag_data[17] = 0;
            rom_imag_data[18] = 0;
            rom_imag_data[19] = 0;
            rom_imag_data[20] = 0;
            rom_imag_data[21] = 0;
            rom_imag_data[22] = 0;
            rom_imag_data[23] = 0;
            rom_imag_data[24] = 0;
            rom_imag_data[25] = 0;
            rom_imag_data[26] = 0;
            rom_imag_data[27] = 0;
            rom_imag_data[28] = 0;
            rom_imag_data[29] = 0;
            rom_imag_data[30] = 0;
            rom_imag_data[31] = 0;
            rom_imag_data[32] = 0;
            rom_imag_data[33] = 0;
            rom_imag_data[34] = 0;
            rom_imag_data[35] = 0;
            rom_imag_data[36] = 0;
            rom_imag_data[37] = 0;
            rom_imag_data[38] = 0;
            rom_imag_data[39] = 0;
            rom_imag_data[40] = 0;
            rom_imag_data[41] = 0;
            rom_imag_data[42] = 0;
            rom_imag_data[43] = 0;
            rom_imag_data[44] = 0;
            rom_imag_data[45] = 0;
            rom_imag_data[46] = 0;
            rom_imag_data[47] = 0;
            rom_imag_data[48] = 0;
            rom_imag_data[49] = 0;
            rom_imag_data[50] = 0;
            rom_imag_data[51] = 0;
            rom_imag_data[52] = 0;
            rom_imag_data[53] = 0;
            rom_imag_data[54] = 0;
            rom_imag_data[55] = 0;
            rom_imag_data[56] = 0;
            rom_imag_data[57] = 0;
            rom_imag_data[58] = 0;
            rom_imag_data[59] = 0;
            rom_imag_data[60] = 0;
            rom_imag_data[61] = 0;
            rom_imag_data[62] = 0;
            rom_imag_data[63] = 0;
            rom_imag_data[64] = 0;
            rom_imag_data[65] = -6;
            rom_imag_data[66] = -13;
            rom_imag_data[67] = -19;
            rom_imag_data[68] = -25;
            rom_imag_data[69] = -31;
            rom_imag_data[70] = -37;
            rom_imag_data[71] = -43;
            rom_imag_data[72] = -49;
            rom_imag_data[73] = -55;
            rom_imag_data[74] = -60;
            rom_imag_data[75] = -66;
            rom_imag_data[76] = -71;
            rom_imag_data[77] = -76;
            rom_imag_data[78] = -81;
            rom_imag_data[79] = -86;
            rom_imag_data[80] = -91;
            rom_imag_data[81] = -95;
            rom_imag_data[82] = -99;
            rom_imag_data[83] = -103;
            rom_imag_data[84] = -106;
            rom_imag_data[85] = -110;
            rom_imag_data[86] = -113;
            rom_imag_data[87] = -116;
            rom_imag_data[88] = -118;
            rom_imag_data[89] = -121;
            rom_imag_data[90] = -122;
            rom_imag_data[91] = -124;
            rom_imag_data[92] = -126;
            rom_imag_data[93] = -127;
            rom_imag_data[94] = -127;
            rom_imag_data[95] = -128;
            rom_imag_data[96] = -128;
            rom_imag_data[97] = -128;
            rom_imag_data[98] = -127;
            rom_imag_data[99] = -127;
            rom_imag_data[100] = -126;
            rom_imag_data[101] = -124;
            rom_imag_data[102] = -122;
            rom_imag_data[103] = -121;
            rom_imag_data[104] = -118;
            rom_imag_data[105] = -116;
            rom_imag_data[106] = -113;
            rom_imag_data[107] = -110;
            rom_imag_data[108] = -106;
            rom_imag_data[109] = -103;
            rom_imag_data[110] = -99;
            rom_imag_data[111] = -95;
            rom_imag_data[112] = -91;
            rom_imag_data[113] = -86;
            rom_imag_data[114] = -81;
            rom_imag_data[115] = -76;
            rom_imag_data[116] = -71;
            rom_imag_data[117] = -66;
            rom_imag_data[118] = -60;
            rom_imag_data[119] = -55;
            rom_imag_data[120] = -49;
            rom_imag_data[121] = -43;
            rom_imag_data[122] = -37;
            rom_imag_data[123] = -31;
            rom_imag_data[124] = -25;
            rom_imag_data[125] = -19;
            rom_imag_data[126] = -13;
            rom_imag_data[127] = -6;
            rom_imag_data[128] = 0;
            rom_imag_data[129] = -3;
            rom_imag_data[130] = -6;
            rom_imag_data[131] = -9;
            rom_imag_data[132] = -13;
            rom_imag_data[133] = -16;
            rom_imag_data[134] = -19;
            rom_imag_data[135] = -22;
            rom_imag_data[136] = -25;
            rom_imag_data[137] = -28;
            rom_imag_data[138] = -31;
            rom_imag_data[139] = -34;
            rom_imag_data[140] = -37;
            rom_imag_data[141] = -40;
            rom_imag_data[142] = -43;
            rom_imag_data[143] = -46;
            rom_imag_data[144] = -49;
            rom_imag_data[145] = -52;
            rom_imag_data[146] = -55;
            rom_imag_data[147] = -58;
            rom_imag_data[148] = -60;
            rom_imag_data[149] = -63;
            rom_imag_data[150] = -66;
            rom_imag_data[151] = -68;
            rom_imag_data[152] = -71;
            rom_imag_data[153] = -74;
            rom_imag_data[154] = -76;
            rom_imag_data[155] = -79;
            rom_imag_data[156] = -81;
            rom_imag_data[157] = -84;
            rom_imag_data[158] = -86;
            rom_imag_data[159] = -88;
            rom_imag_data[160] = -91;
            rom_imag_data[161] = -93;
            rom_imag_data[162] = -95;
            rom_imag_data[163] = -97;
            rom_imag_data[164] = -99;
            rom_imag_data[165] = -101;
            rom_imag_data[166] = -103;
            rom_imag_data[167] = -105;
            rom_imag_data[168] = -106;
            rom_imag_data[169] = -108;
            rom_imag_data[170] = -110;
            rom_imag_data[171] = -111;
            rom_imag_data[172] = -113;
            rom_imag_data[173] = -114;
            rom_imag_data[174] = -116;
            rom_imag_data[175] = -117;
            rom_imag_data[176] = -118;
            rom_imag_data[177] = -119;
            rom_imag_data[178] = -121;
            rom_imag_data[179] = -122;
            rom_imag_data[180] = -122;
            rom_imag_data[181] = -123;
            rom_imag_data[182] = -124;
            rom_imag_data[183] = -125;
            rom_imag_data[184] = -126;
            rom_imag_data[185] = -126;
            rom_imag_data[186] = -127;
            rom_imag_data[187] = -127;
            rom_imag_data[188] = -127;
            rom_imag_data[189] = -128;
            rom_imag_data[190] = -128;
            rom_imag_data[191] = -128;
            rom_imag_data[192] = 0;
            rom_imag_data[193] = -9;
            rom_imag_data[194] = -19;
            rom_imag_data[195] = -28;
            rom_imag_data[196] = -37;
            rom_imag_data[197] = -46;
            rom_imag_data[198] = -55;
            rom_imag_data[199] = -63;
            rom_imag_data[200] = -71;
            rom_imag_data[201] = -79;
            rom_imag_data[202] = -86;
            rom_imag_data[203] = -93;
            rom_imag_data[204] = -99;
            rom_imag_data[205] = -105;
            rom_imag_data[206] = -110;
            rom_imag_data[207] = -114;
            rom_imag_data[208] = -118;
            rom_imag_data[209] = -122;
            rom_imag_data[210] = -124;
            rom_imag_data[211] = -126;
            rom_imag_data[212] = -127;
            rom_imag_data[213] = -128;
            rom_imag_data[214] = -128;
            rom_imag_data[215] = -127;
            rom_imag_data[216] = -126;
            rom_imag_data[217] = -123;
            rom_imag_data[218] = -121;
            rom_imag_data[219] = -117;
            rom_imag_data[220] = -113;
            rom_imag_data[221] = -108;
            rom_imag_data[222] = -103;
            rom_imag_data[223] = -97;
            rom_imag_data[224] = -91;
            rom_imag_data[225] = -84;
            rom_imag_data[226] = -76;
            rom_imag_data[227] = -68;
            rom_imag_data[228] = -60;
            rom_imag_data[229] = -52;
            rom_imag_data[230] = -43;
            rom_imag_data[231] = -34;
            rom_imag_data[232] = -25;
            rom_imag_data[233] = -16;
            rom_imag_data[234] = -6;
            rom_imag_data[235] = 3;
            rom_imag_data[236] = 13;
            rom_imag_data[237] = 22;
            rom_imag_data[238] = 31;
            rom_imag_data[239] = 40;
            rom_imag_data[240] = 49;
            rom_imag_data[241] = 58;
            rom_imag_data[242] = 66;
            rom_imag_data[243] = 74;
            rom_imag_data[244] = 81;
            rom_imag_data[245] = 88;
            rom_imag_data[246] = 95;
            rom_imag_data[247] = 101;
            rom_imag_data[248] = 106;
            rom_imag_data[249] = 111;
            rom_imag_data[250] = 116;
            rom_imag_data[251] = 119;
            rom_imag_data[252] = 122;
            rom_imag_data[253] = 125;
            rom_imag_data[254] = 127;
            rom_imag_data[255] = 128;
            rom_imag_data[256] = 0;
            rom_imag_data[257] = -2;
            rom_imag_data[258] = -3;
            rom_imag_data[259] = -5;
            rom_imag_data[260] = -6;
            rom_imag_data[261] = -8;
            rom_imag_data[262] = -9;
            rom_imag_data[263] = -11;
            rom_imag_data[264] = -13;
            rom_imag_data[265] = -14;
            rom_imag_data[266] = -16;
            rom_imag_data[267] = -17;
            rom_imag_data[268] = -19;
            rom_imag_data[269] = -20;
            rom_imag_data[270] = -22;
            rom_imag_data[271] = -23;
            rom_imag_data[272] = -25;
            rom_imag_data[273] = -27;
            rom_imag_data[274] = -28;
            rom_imag_data[275] = -30;
            rom_imag_data[276] = -31;
            rom_imag_data[277] = -33;
            rom_imag_data[278] = -34;
            rom_imag_data[279] = -36;
            rom_imag_data[280] = -37;
            rom_imag_data[281] = -39;
            rom_imag_data[282] = -40;
            rom_imag_data[283] = -42;
            rom_imag_data[284] = -43;
            rom_imag_data[285] = -45;
            rom_imag_data[286] = -46;
            rom_imag_data[287] = -48;
            rom_imag_data[288] = -49;
            rom_imag_data[289] = -50;
            rom_imag_data[290] = -52;
            rom_imag_data[291] = -53;
            rom_imag_data[292] = -55;
            rom_imag_data[293] = -56;
            rom_imag_data[294] = -58;
            rom_imag_data[295] = -59;
            rom_imag_data[296] = -60;
            rom_imag_data[297] = -62;
            rom_imag_data[298] = -63;
            rom_imag_data[299] = -64;
            rom_imag_data[300] = -66;
            rom_imag_data[301] = -67;
            rom_imag_data[302] = -68;
            rom_imag_data[303] = -70;
            rom_imag_data[304] = -71;
            rom_imag_data[305] = -72;
            rom_imag_data[306] = -74;
            rom_imag_data[307] = -75;
            rom_imag_data[308] = -76;
            rom_imag_data[309] = -78;
            rom_imag_data[310] = -79;
            rom_imag_data[311] = -80;
            rom_imag_data[312] = -81;
            rom_imag_data[313] = -82;
            rom_imag_data[314] = -84;
            rom_imag_data[315] = -85;
            rom_imag_data[316] = -86;
            rom_imag_data[317] = -87;
            rom_imag_data[318] = -88;
            rom_imag_data[319] = -89;
            rom_imag_data[320] = 0;
            rom_imag_data[321] = -8;
            rom_imag_data[322] = -16;
            rom_imag_data[323] = -23;
            rom_imag_data[324] = -31;
            rom_imag_data[325] = -39;
            rom_imag_data[326] = -46;
            rom_imag_data[327] = -53;
            rom_imag_data[328] = -60;
            rom_imag_data[329] = -67;
            rom_imag_data[330] = -74;
            rom_imag_data[331] = -80;
            rom_imag_data[332] = -86;
            rom_imag_data[333] = -92;
            rom_imag_data[334] = -97;
            rom_imag_data[335] = -102;
            rom_imag_data[336] = -106;
            rom_imag_data[337] = -111;
            rom_imag_data[338] = -114;
            rom_imag_data[339] = -118;
            rom_imag_data[340] = -121;
            rom_imag_data[341] = -123;
            rom_imag_data[342] = -125;
            rom_imag_data[343] = -126;
            rom_imag_data[344] = -127;
            rom_imag_data[345] = -128;
            rom_imag_data[346] = -128;
            rom_imag_data[347] = -128;
            rom_imag_data[348] = -127;
            rom_imag_data[349] = -125;
            rom_imag_data[350] = -123;
            rom_imag_data[351] = -121;
            rom_imag_data[352] = -118;
            rom_imag_data[353] = -115;
            rom_imag_data[354] = -111;
            rom_imag_data[355] = -107;
            rom_imag_data[356] = -103;
            rom_imag_data[357] = -98;
            rom_imag_data[358] = -93;
            rom_imag_data[359] = -87;
            rom_imag_data[360] = -81;
            rom_imag_data[361] = -75;
            rom_imag_data[362] = -68;
            rom_imag_data[363] = -62;
            rom_imag_data[364] = -55;
            rom_imag_data[365] = -48;
            rom_imag_data[366] = -40;
            rom_imag_data[367] = -33;
            rom_imag_data[368] = -25;
            rom_imag_data[369] = -17;
            rom_imag_data[370] = -9;
            rom_imag_data[371] = -2;
            rom_imag_data[372] = 6;
            rom_imag_data[373] = 14;
            rom_imag_data[374] = 22;
            rom_imag_data[375] = 30;
            rom_imag_data[376] = 37;
            rom_imag_data[377] = 45;
            rom_imag_data[378] = 52;
            rom_imag_data[379] = 59;
            rom_imag_data[380] = 66;
            rom_imag_data[381] = 72;
            rom_imag_data[382] = 79;
            rom_imag_data[383] = 85;
            rom_imag_data[384] = 0;
            rom_imag_data[385] = -5;
            rom_imag_data[386] = -9;
            rom_imag_data[387] = -14;
            rom_imag_data[388] = -19;
            rom_imag_data[389] = -23;
            rom_imag_data[390] = -28;
            rom_imag_data[391] = -33;
            rom_imag_data[392] = -37;
            rom_imag_data[393] = -42;
            rom_imag_data[394] = -46;
            rom_imag_data[395] = -50;
            rom_imag_data[396] = -55;
            rom_imag_data[397] = -59;
            rom_imag_data[398] = -63;
            rom_imag_data[399] = -67;
            rom_imag_data[400] = -71;
            rom_imag_data[401] = -75;
            rom_imag_data[402] = -79;
            rom_imag_data[403] = -82;
            rom_imag_data[404] = -86;
            rom_imag_data[405] = -89;
            rom_imag_data[406] = -93;
            rom_imag_data[407] = -96;
            rom_imag_data[408] = -99;
            rom_imag_data[409] = -102;
            rom_imag_data[410] = -105;
            rom_imag_data[411] = -107;
            rom_imag_data[412] = -110;
            rom_imag_data[413] = -112;
            rom_imag_data[414] = -114;
            rom_imag_data[415] = -116;
            rom_imag_data[416] = -118;
            rom_imag_data[417] = -120;
            rom_imag_data[418] = -122;
            rom_imag_data[419] = -123;
            rom_imag_data[420] = -124;
            rom_imag_data[421] = -125;
            rom_imag_data[422] = -126;
            rom_imag_data[423] = -127;
            rom_imag_data[424] = -127;
            rom_imag_data[425] = -128;
            rom_imag_data[426] = -128;
            rom_imag_data[427] = -128;
            rom_imag_data[428] = -128;
            rom_imag_data[429] = -128;
            rom_imag_data[430] = -127;
            rom_imag_data[431] = -126;
            rom_imag_data[432] = -126;
            rom_imag_data[433] = -125;
            rom_imag_data[434] = -123;
            rom_imag_data[435] = -122;
            rom_imag_data[436] = -121;
            rom_imag_data[437] = -119;
            rom_imag_data[438] = -117;
            rom_imag_data[439] = -115;
            rom_imag_data[440] = -113;
            rom_imag_data[441] = -111;
            rom_imag_data[442] = -108;
            rom_imag_data[443] = -106;
            rom_imag_data[444] = -103;
            rom_imag_data[445] = -100;
            rom_imag_data[446] = -97;
            rom_imag_data[447] = -94;
            rom_imag_data[448] = 0;
            rom_imag_data[449] = -11;
            rom_imag_data[450] = -22;
            rom_imag_data[451] = -33;
            rom_imag_data[452] = -43;
            rom_imag_data[453] = -53;
            rom_imag_data[454] = -63;
            rom_imag_data[455] = -72;
            rom_imag_data[456] = -81;
            rom_imag_data[457] = -89;
            rom_imag_data[458] = -97;
            rom_imag_data[459] = -104;
            rom_imag_data[460] = -110;
            rom_imag_data[461] = -115;
            rom_imag_data[462] = -119;
            rom_imag_data[463] = -123;
            rom_imag_data[464] = -126;
            rom_imag_data[465] = -127;
            rom_imag_data[466] = -128;
            rom_imag_data[467] = -128;
            rom_imag_data[468] = -127;
            rom_imag_data[469] = -125;
            rom_imag_data[470] = -122;
            rom_imag_data[471] = -118;
            rom_imag_data[472] = -113;
            rom_imag_data[473] = -107;
            rom_imag_data[474] = -101;
            rom_imag_data[475] = -94;
            rom_imag_data[476] = -86;
            rom_imag_data[477] = -78;
            rom_imag_data[478] = -68;
            rom_imag_data[479] = -59;
            rom_imag_data[480] = -49;
            rom_imag_data[481] = -39;
            rom_imag_data[482] = -28;
            rom_imag_data[483] = -17;
            rom_imag_data[484] = -6;
            rom_imag_data[485] = 5;
            rom_imag_data[486] = 16;
            rom_imag_data[487] = 27;
            rom_imag_data[488] = 37;
            rom_imag_data[489] = 48;
            rom_imag_data[490] = 58;
            rom_imag_data[491] = 67;
            rom_imag_data[492] = 76;
            rom_imag_data[493] = 85;
            rom_imag_data[494] = 93;
            rom_imag_data[495] = 100;
            rom_imag_data[496] = 106;
            rom_imag_data[497] = 112;
            rom_imag_data[498] = 117;
            rom_imag_data[499] = 121;
            rom_imag_data[500] = 124;
            rom_imag_data[501] = 126;
            rom_imag_data[502] = 128;
            rom_imag_data[503] = 128;
            rom_imag_data[504] = 127;
            rom_imag_data[505] = 126;
            rom_imag_data[506] = 123;
            rom_imag_data[507] = 120;
            rom_imag_data[508] = 116;
            rom_imag_data[509] = 111;
            rom_imag_data[510] = 105;
            rom_imag_data[511] = 98;
            end
    end

    // always @(posedge clk) begin
    //     twiddle_fac_R_add <= rom_real_data[addr];
    //     twiddle_fac_Q_add <= rom_imag_data[addr];
    //     twiddle_fac_R_sub <= rom_real_data[addr+OFFSET];
    //     twiddle_fac_Q_sub <= rom_imag_data[addr+OFFSET];
    // end

    assign twiddle_fac_R_add = rom_real_data[addr];
    assign twiddle_fac_Q_add = rom_imag_data[addr];
    assign twiddle_fac_R_sub = rom_real_data[addr+OFFSET];
    assign twiddle_fac_Q_sub = rom_imag_data[addr+OFFSET];

endmodule
