`timescale 1ps / 1ps

module rom_twf_gen #(
    parameter ROM_DEPTH = 512,
    parameter TWF_WIDTH = 9,
    parameter ADDR_WIDTH = 9,
    parameter OFFSET = 64
) (
    // input clk,
    input [ADDR_WIDTH-1:0] addr,
    input en,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_R_add,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_Q_add,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_R_sub,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_Q_sub
);

    logic signed [TWF_WIDTH-1:0] rom_real_data[ROM_DEPTH:1];
    logic signed [TWF_WIDTH-1:0] rom_imag_data[ROM_DEPTH:1];

    always @(*) begin
        //initial begin
        if (en) begin
            rom_real_data[1]   = 128;
            rom_real_data[2]   = 128;
            rom_real_data[3]   = 128;
            rom_real_data[4]   = 128;
            rom_real_data[5]   = 128;
            rom_real_data[6]   = 128;
            rom_real_data[7]   = 128;
            rom_real_data[8]   = 128;
            rom_real_data[9]   = 128;
            rom_real_data[10]  = 128;
            rom_real_data[11]  = 128;
            rom_real_data[12]  = 128;
            rom_real_data[13]  = 128;
            rom_real_data[14]  = 128;
            rom_real_data[15]  = 128;
            rom_real_data[16]  = 128;
            rom_real_data[17]  = 128;
            rom_real_data[18]  = 128;
            rom_real_data[19]  = 128;
            rom_real_data[20]  = 128;
            rom_real_data[21]  = 128;
            rom_real_data[22]  = 128;
            rom_real_data[23]  = 128;
            rom_real_data[24]  = 128;
            rom_real_data[25]  = 128;
            rom_real_data[26]  = 128;
            rom_real_data[27]  = 128;
            rom_real_data[28]  = 128;
            rom_real_data[29]  = 128;
            rom_real_data[30]  = 128;
            rom_real_data[31]  = 128;
            rom_real_data[32]  = 128;
            rom_real_data[33]  = 128;
            rom_real_data[34]  = 128;
            rom_real_data[35]  = 128;
            rom_real_data[36]  = 128;
            rom_real_data[37]  = 128;
            rom_real_data[38]  = 128;
            rom_real_data[39]  = 128;
            rom_real_data[40]  = 128;
            rom_real_data[41]  = 128;
            rom_real_data[42]  = 128;
            rom_real_data[43]  = 128;
            rom_real_data[44]  = 128;
            rom_real_data[45]  = 128;
            rom_real_data[46]  = 128;
            rom_real_data[47]  = 128;
            rom_real_data[48]  = 128;
            rom_real_data[49]  = 128;
            rom_real_data[50]  = 128;
            rom_real_data[51]  = 128;
            rom_real_data[52]  = 128;
            rom_real_data[53]  = 128;
            rom_real_data[54]  = 128;
            rom_real_data[55]  = 128;
            rom_real_data[56]  = 128;
            rom_real_data[57]  = 128;
            rom_real_data[58]  = 128;
            rom_real_data[59]  = 128;
            rom_real_data[60]  = 128;
            rom_real_data[61]  = 128;
            rom_real_data[62]  = 128;
            rom_real_data[63]  = 128;
            rom_real_data[64]  = 128;
            rom_real_data[65]  = 128;
            rom_real_data[66]  = 128;
            rom_real_data[67]  = 127;
            rom_real_data[68]  = 127;
            rom_real_data[69]  = 126;
            rom_real_data[70]  = 124;
            rom_real_data[71]  = 122;
            rom_real_data[72]  = 121;
            rom_real_data[73]  = 118;
            rom_real_data[74]  = 116;
            rom_real_data[75]  = 113;
            rom_real_data[76]  = 110;
            rom_real_data[77]  = 106;
            rom_real_data[78]  = 103;
            rom_real_data[79]  = 99;
            rom_real_data[80]  = 95;
            rom_real_data[81]  = 91;
            rom_real_data[82]  = 86;
            rom_real_data[83]  = 81;
            rom_real_data[84]  = 76;
            rom_real_data[85]  = 71;
            rom_real_data[86]  = 66;
            rom_real_data[87]  = 60;
            rom_real_data[88]  = 55;
            rom_real_data[89]  = 49;
            rom_real_data[90]  = 43;
            rom_real_data[91]  = 37;
            rom_real_data[92]  = 31;
            rom_real_data[93]  = 25;
            rom_real_data[94]  = 19;
            rom_real_data[95]  = 13;
            rom_real_data[96]  = 6;
            rom_real_data[97]  = 0;
            rom_real_data[98]  = -6;
            rom_real_data[99]  = -13;
            rom_real_data[100] = -19;
            rom_real_data[101] = -25;
            rom_real_data[102] = -31;
            rom_real_data[103] = -37;
            rom_real_data[104] = -43;
            rom_real_data[105] = -49;
            rom_real_data[106] = -55;
            rom_real_data[107] = -60;
            rom_real_data[108] = -66;
            rom_real_data[109] = -71;
            rom_real_data[110] = -76;
            rom_real_data[111] = -81;
            rom_real_data[112] = -86;
            rom_real_data[113] = -91;
            rom_real_data[114] = -95;
            rom_real_data[115] = -99;
            rom_real_data[116] = -103;
            rom_real_data[117] = -106;
            rom_real_data[118] = -110;
            rom_real_data[119] = -113;
            rom_real_data[120] = -116;
            rom_real_data[121] = -118;
            rom_real_data[122] = -121;
            rom_real_data[123] = -122;
            rom_real_data[124] = -124;
            rom_real_data[125] = -126;
            rom_real_data[126] = -127;
            rom_real_data[127] = -127;
            rom_real_data[128] = -128;
            rom_real_data[129] = 128;
            rom_real_data[130] = 128;
            rom_real_data[131] = 128;
            rom_real_data[132] = 128;
            rom_real_data[133] = 127;
            rom_real_data[134] = 127;
            rom_real_data[135] = 127;
            rom_real_data[136] = 126;
            rom_real_data[137] = 126;
            rom_real_data[138] = 125;
            rom_real_data[139] = 124;
            rom_real_data[140] = 123;
            rom_real_data[141] = 122;
            rom_real_data[142] = 122;
            rom_real_data[143] = 121;
            rom_real_data[144] = 119;
            rom_real_data[145] = 118;
            rom_real_data[146] = 117;
            rom_real_data[147] = 116;
            rom_real_data[148] = 114;
            rom_real_data[149] = 113;
            rom_real_data[150] = 111;
            rom_real_data[151] = 110;
            rom_real_data[152] = 108;
            rom_real_data[153] = 106;
            rom_real_data[154] = 105;
            rom_real_data[155] = 103;
            rom_real_data[156] = 101;
            rom_real_data[157] = 99;
            rom_real_data[158] = 97;
            rom_real_data[159] = 95;
            rom_real_data[160] = 93;
            rom_real_data[161] = 91;
            rom_real_data[162] = 88;
            rom_real_data[163] = 86;
            rom_real_data[164] = 84;
            rom_real_data[165] = 81;
            rom_real_data[166] = 79;
            rom_real_data[167] = 76;
            rom_real_data[168] = 74;
            rom_real_data[169] = 71;
            rom_real_data[170] = 68;
            rom_real_data[171] = 66;
            rom_real_data[172] = 63;
            rom_real_data[173] = 60;
            rom_real_data[174] = 58;
            rom_real_data[175] = 55;
            rom_real_data[176] = 52;
            rom_real_data[177] = 49;
            rom_real_data[178] = 46;
            rom_real_data[179] = 43;
            rom_real_data[180] = 40;
            rom_real_data[181] = 37;
            rom_real_data[182] = 34;
            rom_real_data[183] = 31;
            rom_real_data[184] = 28;
            rom_real_data[185] = 25;
            rom_real_data[186] = 22;
            rom_real_data[187] = 19;
            rom_real_data[188] = 16;
            rom_real_data[189] = 13;
            rom_real_data[190] = 9;
            rom_real_data[191] = 6;
            rom_real_data[192] = 3;
            rom_real_data[193] = 128;
            rom_real_data[194] = 128;
            rom_real_data[195] = 127;
            rom_real_data[196] = 125;
            rom_real_data[197] = 122;
            rom_real_data[198] = 119;
            rom_real_data[199] = 116;
            rom_real_data[200] = 111;
            rom_real_data[201] = 106;
            rom_real_data[202] = 101;
            rom_real_data[203] = 95;
            rom_real_data[204] = 88;
            rom_real_data[205] = 81;
            rom_real_data[206] = 74;
            rom_real_data[207] = 66;
            rom_real_data[208] = 58;
            rom_real_data[209] = 49;
            rom_real_data[210] = 40;
            rom_real_data[211] = 31;
            rom_real_data[212] = 22;
            rom_real_data[213] = 13;
            rom_real_data[214] = 3;
            rom_real_data[215] = -6;
            rom_real_data[216] = -16;
            rom_real_data[217] = -25;
            rom_real_data[218] = -34;
            rom_real_data[219] = -43;
            rom_real_data[220] = -52;
            rom_real_data[221] = -60;
            rom_real_data[222] = -68;
            rom_real_data[223] = -76;
            rom_real_data[224] = -84;
            rom_real_data[225] = -91;
            rom_real_data[226] = -97;
            rom_real_data[227] = -103;
            rom_real_data[228] = -108;
            rom_real_data[229] = -113;
            rom_real_data[230] = -117;
            rom_real_data[231] = -121;
            rom_real_data[232] = -123;
            rom_real_data[233] = -126;
            rom_real_data[234] = -127;
            rom_real_data[235] = -128;
            rom_real_data[236] = -128;
            rom_real_data[237] = -127;
            rom_real_data[238] = -126;
            rom_real_data[239] = -124;
            rom_real_data[240] = -122;
            rom_real_data[241] = -118;
            rom_real_data[242] = -114;
            rom_real_data[243] = -110;
            rom_real_data[244] = -105;
            rom_real_data[245] = -99;
            rom_real_data[246] = -93;
            rom_real_data[247] = -86;
            rom_real_data[248] = -79;
            rom_real_data[249] = -71;
            rom_real_data[250] = -63;
            rom_real_data[251] = -55;
            rom_real_data[252] = -46;
            rom_real_data[253] = -37;
            rom_real_data[254] = -28;
            rom_real_data[255] = -19;
            rom_real_data[256] = -9;
            rom_real_data[257] = 128;
            rom_real_data[258] = 128;
            rom_real_data[259] = 128;
            rom_real_data[260] = 128;
            rom_real_data[261] = 128;
            rom_real_data[262] = 128;
            rom_real_data[263] = 128;
            rom_real_data[264] = 128;
            rom_real_data[265] = 127;
            rom_real_data[266] = 127;
            rom_real_data[267] = 127;
            rom_real_data[268] = 127;
            rom_real_data[269] = 127;
            rom_real_data[270] = 126;
            rom_real_data[271] = 126;
            rom_real_data[272] = 126;
            rom_real_data[273] = 126;
            rom_real_data[274] = 125;
            rom_real_data[275] = 125;
            rom_real_data[276] = 125;
            rom_real_data[277] = 124;
            rom_real_data[278] = 124;
            rom_real_data[279] = 123;
            rom_real_data[280] = 123;
            rom_real_data[281] = 122;
            rom_real_data[282] = 122;
            rom_real_data[283] = 122;
            rom_real_data[284] = 121;
            rom_real_data[285] = 121;
            rom_real_data[286] = 120;
            rom_real_data[287] = 119;
            rom_real_data[288] = 119;
            rom_real_data[289] = 118;
            rom_real_data[290] = 118;
            rom_real_data[291] = 117;
            rom_real_data[292] = 116;
            rom_real_data[293] = 116;
            rom_real_data[294] = 115;
            rom_real_data[295] = 114;
            rom_real_data[296] = 114;
            rom_real_data[297] = 113;
            rom_real_data[298] = 112;
            rom_real_data[299] = 111;
            rom_real_data[300] = 111;
            rom_real_data[301] = 110;
            rom_real_data[302] = 109;
            rom_real_data[303] = 108;
            rom_real_data[304] = 107;
            rom_real_data[305] = 106;
            rom_real_data[306] = 106;
            rom_real_data[307] = 105;
            rom_real_data[308] = 104;
            rom_real_data[309] = 103;
            rom_real_data[310] = 102;
            rom_real_data[311] = 101;
            rom_real_data[312] = 100;
            rom_real_data[313] = 99;
            rom_real_data[314] = 98;
            rom_real_data[315] = 97;
            rom_real_data[316] = 96;
            rom_real_data[317] = 95;
            rom_real_data[318] = 94;
            rom_real_data[319] = 93;
            rom_real_data[320] = 92;
            rom_real_data[321] = 128;
            rom_real_data[322] = 128;
            rom_real_data[323] = 127;
            rom_real_data[324] = 126;
            rom_real_data[325] = 124;
            rom_real_data[326] = 122;
            rom_real_data[327] = 119;
            rom_real_data[328] = 116;
            rom_real_data[329] = 113;
            rom_real_data[330] = 109;
            rom_real_data[331] = 105;
            rom_real_data[332] = 100;
            rom_real_data[333] = 95;
            rom_real_data[334] = 89;
            rom_real_data[335] = 84;
            rom_real_data[336] = 78;
            rom_real_data[337] = 71;
            rom_real_data[338] = 64;
            rom_real_data[339] = 58;
            rom_real_data[340] = 50;
            rom_real_data[341] = 43;
            rom_real_data[342] = 36;
            rom_real_data[343] = 28;
            rom_real_data[344] = 20;
            rom_real_data[345] = 13;
            rom_real_data[346] = 5;
            rom_real_data[347] = -3;
            rom_real_data[348] = -11;
            rom_real_data[349] = -19;
            rom_real_data[350] = -27;
            rom_real_data[351] = -34;
            rom_real_data[352] = -42;
            rom_real_data[353] = -49;
            rom_real_data[354] = -56;
            rom_real_data[355] = -63;
            rom_real_data[356] = -70;
            rom_real_data[357] = -76;
            rom_real_data[358] = -82;
            rom_real_data[359] = -88;
            rom_real_data[360] = -94;
            rom_real_data[361] = -99;
            rom_real_data[362] = -104;
            rom_real_data[363] = -108;
            rom_real_data[364] = -112;
            rom_real_data[365] = -116;
            rom_real_data[366] = -119;
            rom_real_data[367] = -122;
            rom_real_data[368] = -124;
            rom_real_data[369] = -126;
            rom_real_data[370] = -127;
            rom_real_data[371] = -128;
            rom_real_data[372] = -128;
            rom_real_data[373] = -128;
            rom_real_data[374] = -127;
            rom_real_data[375] = -126;
            rom_real_data[376] = -125;
            rom_real_data[377] = -122;
            rom_real_data[378] = -120;
            rom_real_data[379] = -117;
            rom_real_data[380] = -114;
            rom_real_data[381] = -110;
            rom_real_data[382] = -106;
            rom_real_data[383] = -101;
            rom_real_data[384] = -96;
            rom_real_data[385] = 128;
            rom_real_data[386] = 128;
            rom_real_data[387] = 128;
            rom_real_data[388] = 127;
            rom_real_data[389] = 127;
            rom_real_data[390] = 126;
            rom_real_data[391] = 125;
            rom_real_data[392] = 124;
            rom_real_data[393] = 122;
            rom_real_data[394] = 121;
            rom_real_data[395] = 119;
            rom_real_data[396] = 118;
            rom_real_data[397] = 116;
            rom_real_data[398] = 114;
            rom_real_data[399] = 111;
            rom_real_data[400] = 109;
            rom_real_data[401] = 106;
            rom_real_data[402] = 104;
            rom_real_data[403] = 101;
            rom_real_data[404] = 98;
            rom_real_data[405] = 95;
            rom_real_data[406] = 92;
            rom_real_data[407] = 88;
            rom_real_data[408] = 85;
            rom_real_data[409] = 81;
            rom_real_data[410] = 78;
            rom_real_data[411] = 74;
            rom_real_data[412] = 70;
            rom_real_data[413] = 66;
            rom_real_data[414] = 62;
            rom_real_data[415] = 58;
            rom_real_data[416] = 53;
            rom_real_data[417] = 49;
            rom_real_data[418] = 45;
            rom_real_data[419] = 40;
            rom_real_data[420] = 36;
            rom_real_data[421] = 31;
            rom_real_data[422] = 27;
            rom_real_data[423] = 22;
            rom_real_data[424] = 17;
            rom_real_data[425] = 13;
            rom_real_data[426] = 8;
            rom_real_data[427] = 3;
            rom_real_data[428] = -2;
            rom_real_data[429] = -6;
            rom_real_data[430] = -11;
            rom_real_data[431] = -16;
            rom_real_data[432] = -20;
            rom_real_data[433] = -25;
            rom_real_data[434] = -30;
            rom_real_data[435] = -34;
            rom_real_data[436] = -39;
            rom_real_data[437] = -43;
            rom_real_data[438] = -48;
            rom_real_data[439] = -52;
            rom_real_data[440] = -56;
            rom_real_data[441] = -60;
            rom_real_data[442] = -64;
            rom_real_data[443] = -68;
            rom_real_data[444] = -72;
            rom_real_data[445] = -76;
            rom_real_data[446] = -80;
            rom_real_data[447] = -84;
            rom_real_data[448] = -87;
            rom_real_data[449] = 128;
            rom_real_data[450] = 128;
            rom_real_data[451] = 126;
            rom_real_data[452] = 124;
            rom_real_data[453] = 121;
            rom_real_data[454] = 116;
            rom_real_data[455] = 111;
            rom_real_data[456] = 106;
            rom_real_data[457] = 99;
            rom_real_data[458] = 92;
            rom_real_data[459] = 84;
            rom_real_data[460] = 75;
            rom_real_data[461] = 66;
            rom_real_data[462] = 56;
            rom_real_data[463] = 46;
            rom_real_data[464] = 36;
            rom_real_data[465] = 25;
            rom_real_data[466] = 14;
            rom_real_data[467] = 3;
            rom_real_data[468] = -8;
            rom_real_data[469] = -19;
            rom_real_data[470] = -30;
            rom_real_data[471] = -40;
            rom_real_data[472] = -50;
            rom_real_data[473] = -60;
            rom_real_data[474] = -70;
            rom_real_data[475] = -79;
            rom_real_data[476] = -87;
            rom_real_data[477] = -95;
            rom_real_data[478] = -102;
            rom_real_data[479] = -108;
            rom_real_data[480] = -114;
            rom_real_data[481] = -118;
            rom_real_data[482] = -122;
            rom_real_data[483] = -125;
            rom_real_data[484] = -127;
            rom_real_data[485] = -128;
            rom_real_data[486] = -128;
            rom_real_data[487] = -127;
            rom_real_data[488] = -125;
            rom_real_data[489] = -122;
            rom_real_data[490] = -119;
            rom_real_data[491] = -114;
            rom_real_data[492] = -109;
            rom_real_data[493] = -103;
            rom_real_data[494] = -96;
            rom_real_data[495] = -88;
            rom_real_data[496] = -80;
            rom_real_data[497] = -71;
            rom_real_data[498] = -62;
            rom_real_data[499] = -52;
            rom_real_data[500] = -42;
            rom_real_data[501] = -31;
            rom_real_data[502] = -20;
            rom_real_data[503] = -9;
            rom_real_data[504] = 2;
            rom_real_data[505] = 13;
            rom_real_data[506] = 23;
            rom_real_data[507] = 34;
            rom_real_data[508] = 45;
            rom_real_data[509] = 55;
            rom_real_data[510] = 64;
            rom_real_data[511] = 74;
            rom_real_data[512] = 82;


            rom_imag_data[1]   = 0;
            rom_imag_data[2]   = 0;
            rom_imag_data[3]   = 0;
            rom_imag_data[4]   = 0;
            rom_imag_data[5]   = 0;
            rom_imag_data[6]   = 0;
            rom_imag_data[7]   = 0;
            rom_imag_data[8]   = 0;
            rom_imag_data[9]   = 0;
            rom_imag_data[10]  = 0;
            rom_imag_data[11]  = 0;
            rom_imag_data[12]  = 0;
            rom_imag_data[13]  = 0;
            rom_imag_data[14]  = 0;
            rom_imag_data[15]  = 0;
            rom_imag_data[16]  = 0;
            rom_imag_data[17]  = 0;
            rom_imag_data[18]  = 0;
            rom_imag_data[19]  = 0;
            rom_imag_data[20]  = 0;
            rom_imag_data[21]  = 0;
            rom_imag_data[22]  = 0;
            rom_imag_data[23]  = 0;
            rom_imag_data[24]  = 0;
            rom_imag_data[25]  = 0;
            rom_imag_data[26]  = 0;
            rom_imag_data[27]  = 0;
            rom_imag_data[28]  = 0;
            rom_imag_data[29]  = 0;
            rom_imag_data[30]  = 0;
            rom_imag_data[31]  = 0;
            rom_imag_data[32]  = 0;
            rom_imag_data[33]  = 0;
            rom_imag_data[34]  = 0;
            rom_imag_data[35]  = 0;
            rom_imag_data[36]  = 0;
            rom_imag_data[37]  = 0;
            rom_imag_data[38]  = 0;
            rom_imag_data[39]  = 0;
            rom_imag_data[40]  = 0;
            rom_imag_data[41]  = 0;
            rom_imag_data[42]  = 0;
            rom_imag_data[43]  = 0;
            rom_imag_data[44]  = 0;
            rom_imag_data[45]  = 0;
            rom_imag_data[46]  = 0;
            rom_imag_data[47]  = 0;
            rom_imag_data[48]  = 0;
            rom_imag_data[49]  = 0;
            rom_imag_data[50]  = 0;
            rom_imag_data[51]  = 0;
            rom_imag_data[52]  = 0;
            rom_imag_data[53]  = 0;
            rom_imag_data[54]  = 0;
            rom_imag_data[55]  = 0;
            rom_imag_data[56]  = 0;
            rom_imag_data[57]  = 0;
            rom_imag_data[58]  = 0;
            rom_imag_data[59]  = 0;
            rom_imag_data[60]  = 0;
            rom_imag_data[61]  = 0;
            rom_imag_data[62]  = 0;
            rom_imag_data[63]  = 0;
            rom_imag_data[64]  = 0;
            rom_imag_data[65]  = 0;
            rom_imag_data[66]  = -6;
            rom_imag_data[67]  = -13;
            rom_imag_data[68]  = -19;
            rom_imag_data[69]  = -25;
            rom_imag_data[70]  = -31;
            rom_imag_data[71]  = -37;
            rom_imag_data[72]  = -43;
            rom_imag_data[73]  = -49;
            rom_imag_data[74]  = -55;
            rom_imag_data[75]  = -60;
            rom_imag_data[76]  = -66;
            rom_imag_data[77]  = -71;
            rom_imag_data[78]  = -76;
            rom_imag_data[79]  = -81;
            rom_imag_data[80]  = -86;
            rom_imag_data[81]  = -91;
            rom_imag_data[82]  = -95;
            rom_imag_data[83]  = -99;
            rom_imag_data[84]  = -103;
            rom_imag_data[85]  = -106;
            rom_imag_data[86]  = -110;
            rom_imag_data[87]  = -113;
            rom_imag_data[88]  = -116;
            rom_imag_data[89]  = -118;
            rom_imag_data[90]  = -121;
            rom_imag_data[91]  = -122;
            rom_imag_data[92]  = -124;
            rom_imag_data[93]  = -126;
            rom_imag_data[94]  = -127;
            rom_imag_data[95]  = -127;
            rom_imag_data[96]  = -128;
            rom_imag_data[97]  = -128;
            rom_imag_data[98]  = -128;
            rom_imag_data[99]  = -127;
            rom_imag_data[100] = -127;
            rom_imag_data[101] = -126;
            rom_imag_data[102] = -124;
            rom_imag_data[103] = -122;
            rom_imag_data[104] = -121;
            rom_imag_data[105] = -118;
            rom_imag_data[106] = -116;
            rom_imag_data[107] = -113;
            rom_imag_data[108] = -110;
            rom_imag_data[109] = -106;
            rom_imag_data[110] = -103;
            rom_imag_data[111] = -99;
            rom_imag_data[112] = -95;
            rom_imag_data[113] = -91;
            rom_imag_data[114] = -86;
            rom_imag_data[115] = -81;
            rom_imag_data[116] = -76;
            rom_imag_data[117] = -71;
            rom_imag_data[118] = -66;
            rom_imag_data[119] = -60;
            rom_imag_data[120] = -55;
            rom_imag_data[121] = -49;
            rom_imag_data[122] = -43;
            rom_imag_data[123] = -37;
            rom_imag_data[124] = -31;
            rom_imag_data[125] = -25;
            rom_imag_data[126] = -19;
            rom_imag_data[127] = -13;
            rom_imag_data[128] = -6;
            rom_imag_data[129] = 0;
            rom_imag_data[130] = -3;
            rom_imag_data[131] = -6;
            rom_imag_data[132] = -9;
            rom_imag_data[133] = -13;
            rom_imag_data[134] = -16;
            rom_imag_data[135] = -19;
            rom_imag_data[136] = -22;
            rom_imag_data[137] = -25;
            rom_imag_data[138] = -28;
            rom_imag_data[139] = -31;
            rom_imag_data[140] = -34;
            rom_imag_data[141] = -37;
            rom_imag_data[142] = -40;
            rom_imag_data[143] = -43;
            rom_imag_data[144] = -46;
            rom_imag_data[145] = -49;
            rom_imag_data[146] = -52;
            rom_imag_data[147] = -55;
            rom_imag_data[148] = -58;
            rom_imag_data[149] = -60;
            rom_imag_data[150] = -63;
            rom_imag_data[151] = -66;
            rom_imag_data[152] = -68;
            rom_imag_data[153] = -71;
            rom_imag_data[154] = -74;
            rom_imag_data[155] = -76;
            rom_imag_data[156] = -79;
            rom_imag_data[157] = -81;
            rom_imag_data[158] = -84;
            rom_imag_data[159] = -86;
            rom_imag_data[160] = -88;
            rom_imag_data[161] = -91;
            rom_imag_data[162] = -93;
            rom_imag_data[163] = -95;
            rom_imag_data[164] = -97;
            rom_imag_data[165] = -99;
            rom_imag_data[166] = -101;
            rom_imag_data[167] = -103;
            rom_imag_data[168] = -105;
            rom_imag_data[169] = -106;
            rom_imag_data[170] = -108;
            rom_imag_data[171] = -110;
            rom_imag_data[172] = -111;
            rom_imag_data[173] = -113;
            rom_imag_data[174] = -114;
            rom_imag_data[175] = -116;
            rom_imag_data[176] = -117;
            rom_imag_data[177] = -118;
            rom_imag_data[178] = -119;
            rom_imag_data[179] = -121;
            rom_imag_data[180] = -122;
            rom_imag_data[181] = -122;
            rom_imag_data[182] = -123;
            rom_imag_data[183] = -124;
            rom_imag_data[184] = -125;
            rom_imag_data[185] = -126;
            rom_imag_data[186] = -126;
            rom_imag_data[187] = -127;
            rom_imag_data[188] = -127;
            rom_imag_data[189] = -127;
            rom_imag_data[190] = -128;
            rom_imag_data[191] = -128;
            rom_imag_data[192] = -128;
            rom_imag_data[193] = 0;
            rom_imag_data[194] = -9;
            rom_imag_data[195] = -19;
            rom_imag_data[196] = -28;
            rom_imag_data[197] = -37;
            rom_imag_data[198] = -46;
            rom_imag_data[199] = -55;
            rom_imag_data[200] = -63;
            rom_imag_data[201] = -71;
            rom_imag_data[202] = -79;
            rom_imag_data[203] = -86;
            rom_imag_data[204] = -93;
            rom_imag_data[205] = -99;
            rom_imag_data[206] = -105;
            rom_imag_data[207] = -110;
            rom_imag_data[208] = -114;
            rom_imag_data[209] = -118;
            rom_imag_data[210] = -122;
            rom_imag_data[211] = -124;
            rom_imag_data[212] = -126;
            rom_imag_data[213] = -127;
            rom_imag_data[214] = -128;
            rom_imag_data[215] = -128;
            rom_imag_data[216] = -127;
            rom_imag_data[217] = -126;
            rom_imag_data[218] = -123;
            rom_imag_data[219] = -121;
            rom_imag_data[220] = -117;
            rom_imag_data[221] = -113;
            rom_imag_data[222] = -108;
            rom_imag_data[223] = -103;
            rom_imag_data[224] = -97;
            rom_imag_data[225] = -91;
            rom_imag_data[226] = -84;
            rom_imag_data[227] = -76;
            rom_imag_data[228] = -68;
            rom_imag_data[229] = -60;
            rom_imag_data[230] = -52;
            rom_imag_data[231] = -43;
            rom_imag_data[232] = -34;
            rom_imag_data[233] = -25;
            rom_imag_data[234] = -16;
            rom_imag_data[235] = -6;
            rom_imag_data[236] = 3;
            rom_imag_data[237] = 13;
            rom_imag_data[238] = 22;
            rom_imag_data[239] = 31;
            rom_imag_data[240] = 40;
            rom_imag_data[241] = 49;
            rom_imag_data[242] = 58;
            rom_imag_data[243] = 66;
            rom_imag_data[244] = 74;
            rom_imag_data[245] = 81;
            rom_imag_data[246] = 88;
            rom_imag_data[247] = 95;
            rom_imag_data[248] = 101;
            rom_imag_data[249] = 106;
            rom_imag_data[250] = 111;
            rom_imag_data[251] = 116;
            rom_imag_data[252] = 119;
            rom_imag_data[253] = 122;
            rom_imag_data[254] = 125;
            rom_imag_data[255] = 127;
            rom_imag_data[256] = 128;
            rom_imag_data[257] = 0;
            rom_imag_data[258] = -2;
            rom_imag_data[259] = -3;
            rom_imag_data[260] = -5;
            rom_imag_data[261] = -6;
            rom_imag_data[262] = -8;
            rom_imag_data[263] = -9;
            rom_imag_data[264] = -11;
            rom_imag_data[265] = -13;
            rom_imag_data[266] = -14;
            rom_imag_data[267] = -16;
            rom_imag_data[268] = -17;
            rom_imag_data[269] = -19;
            rom_imag_data[270] = -20;
            rom_imag_data[271] = -22;
            rom_imag_data[272] = -23;
            rom_imag_data[273] = -25;
            rom_imag_data[274] = -27;
            rom_imag_data[275] = -28;
            rom_imag_data[276] = -30;
            rom_imag_data[277] = -31;
            rom_imag_data[278] = -33;
            rom_imag_data[279] = -34;
            rom_imag_data[280] = -36;
            rom_imag_data[281] = -37;
            rom_imag_data[282] = -39;
            rom_imag_data[283] = -40;
            rom_imag_data[284] = -42;
            rom_imag_data[285] = -43;
            rom_imag_data[286] = -45;
            rom_imag_data[287] = -46;
            rom_imag_data[288] = -48;
            rom_imag_data[289] = -49;
            rom_imag_data[290] = -50;
            rom_imag_data[291] = -52;
            rom_imag_data[292] = -53;
            rom_imag_data[293] = -55;
            rom_imag_data[294] = -56;
            rom_imag_data[295] = -58;
            rom_imag_data[296] = -59;
            rom_imag_data[297] = -60;
            rom_imag_data[298] = -62;
            rom_imag_data[299] = -63;
            rom_imag_data[300] = -64;
            rom_imag_data[301] = -66;
            rom_imag_data[302] = -67;
            rom_imag_data[303] = -68;
            rom_imag_data[304] = -70;
            rom_imag_data[305] = -71;
            rom_imag_data[306] = -72;
            rom_imag_data[307] = -74;
            rom_imag_data[308] = -75;
            rom_imag_data[309] = -76;
            rom_imag_data[310] = -78;
            rom_imag_data[311] = -79;
            rom_imag_data[312] = -80;
            rom_imag_data[313] = -81;
            rom_imag_data[314] = -82;
            rom_imag_data[315] = -84;
            rom_imag_data[316] = -85;
            rom_imag_data[317] = -86;
            rom_imag_data[318] = -87;
            rom_imag_data[319] = -88;
            rom_imag_data[320] = -89;
            rom_imag_data[321] = 0;
            rom_imag_data[322] = -8;
            rom_imag_data[323] = -16;
            rom_imag_data[324] = -23;
            rom_imag_data[325] = -31;
            rom_imag_data[326] = -39;
            rom_imag_data[327] = -46;
            rom_imag_data[328] = -53;
            rom_imag_data[329] = -60;
            rom_imag_data[330] = -67;
            rom_imag_data[331] = -74;
            rom_imag_data[332] = -80;
            rom_imag_data[333] = -86;
            rom_imag_data[334] = -92;
            rom_imag_data[335] = -97;
            rom_imag_data[336] = -102;
            rom_imag_data[337] = -106;
            rom_imag_data[338] = -111;
            rom_imag_data[339] = -114;
            rom_imag_data[340] = -118;
            rom_imag_data[341] = -121;
            rom_imag_data[342] = -123;
            rom_imag_data[343] = -125;
            rom_imag_data[344] = -126;
            rom_imag_data[345] = -127;
            rom_imag_data[346] = -128;
            rom_imag_data[347] = -128;
            rom_imag_data[348] = -128;
            rom_imag_data[349] = -127;
            rom_imag_data[350] = -125;
            rom_imag_data[351] = -123;
            rom_imag_data[352] = -121;
            rom_imag_data[353] = -118;
            rom_imag_data[354] = -115;
            rom_imag_data[355] = -111;
            rom_imag_data[356] = -107;
            rom_imag_data[357] = -103;
            rom_imag_data[358] = -98;
            rom_imag_data[359] = -93;
            rom_imag_data[360] = -87;
            rom_imag_data[361] = -81;
            rom_imag_data[362] = -75;
            rom_imag_data[363] = -68;
            rom_imag_data[364] = -62;
            rom_imag_data[365] = -55;
            rom_imag_data[366] = -48;
            rom_imag_data[367] = -40;
            rom_imag_data[368] = -33;
            rom_imag_data[369] = -25;
            rom_imag_data[370] = -17;
            rom_imag_data[371] = -9;
            rom_imag_data[372] = -2;
            rom_imag_data[373] = 6;
            rom_imag_data[374] = 14;
            rom_imag_data[375] = 22;
            rom_imag_data[376] = 30;
            rom_imag_data[377] = 37;
            rom_imag_data[378] = 45;
            rom_imag_data[379] = 52;
            rom_imag_data[380] = 59;
            rom_imag_data[381] = 66;
            rom_imag_data[382] = 72;
            rom_imag_data[383] = 79;
            rom_imag_data[384] = 85;
            rom_imag_data[385] = 0;
            rom_imag_data[386] = -5;
            rom_imag_data[387] = -9;
            rom_imag_data[388] = -14;
            rom_imag_data[389] = -19;
            rom_imag_data[390] = -23;
            rom_imag_data[391] = -28;
            rom_imag_data[392] = -33;
            rom_imag_data[393] = -37;
            rom_imag_data[394] = -42;
            rom_imag_data[395] = -46;
            rom_imag_data[396] = -50;
            rom_imag_data[397] = -55;
            rom_imag_data[398] = -59;
            rom_imag_data[399] = -63;
            rom_imag_data[400] = -67;
            rom_imag_data[401] = -71;
            rom_imag_data[402] = -75;
            rom_imag_data[403] = -79;
            rom_imag_data[404] = -82;
            rom_imag_data[405] = -86;
            rom_imag_data[406] = -89;
            rom_imag_data[407] = -93;
            rom_imag_data[408] = -96;
            rom_imag_data[409] = -99;
            rom_imag_data[410] = -102;
            rom_imag_data[411] = -105;
            rom_imag_data[412] = -107;
            rom_imag_data[413] = -110;
            rom_imag_data[414] = -112;
            rom_imag_data[415] = -114;
            rom_imag_data[416] = -116;
            rom_imag_data[417] = -118;
            rom_imag_data[418] = -120;
            rom_imag_data[419] = -122;
            rom_imag_data[420] = -123;
            rom_imag_data[421] = -124;
            rom_imag_data[422] = -125;
            rom_imag_data[423] = -126;
            rom_imag_data[424] = -127;
            rom_imag_data[425] = -127;
            rom_imag_data[426] = -128;
            rom_imag_data[427] = -128;
            rom_imag_data[428] = -128;
            rom_imag_data[429] = -128;
            rom_imag_data[430] = -128;
            rom_imag_data[431] = -127;
            rom_imag_data[432] = -126;
            rom_imag_data[433] = -126;
            rom_imag_data[434] = -125;
            rom_imag_data[435] = -123;
            rom_imag_data[436] = -122;
            rom_imag_data[437] = -121;
            rom_imag_data[438] = -119;
            rom_imag_data[439] = -117;
            rom_imag_data[440] = -115;
            rom_imag_data[441] = -113;
            rom_imag_data[442] = -111;
            rom_imag_data[443] = -108;
            rom_imag_data[444] = -106;
            rom_imag_data[445] = -103;
            rom_imag_data[446] = -100;
            rom_imag_data[447] = -97;
            rom_imag_data[448] = -94;
            rom_imag_data[449] = 0;
            rom_imag_data[450] = -11;
            rom_imag_data[451] = -22;
            rom_imag_data[452] = -33;
            rom_imag_data[453] = -43;
            rom_imag_data[454] = -53;
            rom_imag_data[455] = -63;
            rom_imag_data[456] = -72;
            rom_imag_data[457] = -81;
            rom_imag_data[458] = -89;
            rom_imag_data[459] = -97;
            rom_imag_data[460] = -104;
            rom_imag_data[461] = -110;
            rom_imag_data[462] = -115;
            rom_imag_data[463] = -119;
            rom_imag_data[464] = -123;
            rom_imag_data[465] = -126;
            rom_imag_data[466] = -127;
            rom_imag_data[467] = -128;
            rom_imag_data[468] = -128;
            rom_imag_data[469] = -127;
            rom_imag_data[470] = -125;
            rom_imag_data[471] = -122;
            rom_imag_data[472] = -118;
            rom_imag_data[473] = -113;
            rom_imag_data[474] = -107;
            rom_imag_data[475] = -101;
            rom_imag_data[476] = -94;
            rom_imag_data[477] = -86;
            rom_imag_data[478] = -78;
            rom_imag_data[479] = -68;
            rom_imag_data[480] = -59;
            rom_imag_data[481] = -49;
            rom_imag_data[482] = -39;
            rom_imag_data[483] = -28;
            rom_imag_data[484] = -17;
            rom_imag_data[485] = -6;
            rom_imag_data[486] = 5;
            rom_imag_data[487] = 16;
            rom_imag_data[488] = 27;
            rom_imag_data[489] = 37;
            rom_imag_data[490] = 48;
            rom_imag_data[491] = 58;
            rom_imag_data[492] = 67;
            rom_imag_data[493] = 76;
            rom_imag_data[494] = 85;
            rom_imag_data[495] = 93;
            rom_imag_data[496] = 100;
            rom_imag_data[497] = 106;
            rom_imag_data[498] = 112;
            rom_imag_data[499] = 117;
            rom_imag_data[500] = 121;
            rom_imag_data[501] = 124;
            rom_imag_data[502] = 126;
            rom_imag_data[503] = 128;
            rom_imag_data[504] = 128;
            rom_imag_data[505] = 127;
            rom_imag_data[506] = 126;
            rom_imag_data[507] = 123;
            rom_imag_data[508] = 120;
            rom_imag_data[509] = 116;
            rom_imag_data[510] = 111;
            rom_imag_data[511] = 105;
            rom_imag_data[512] = 98;
        end
    end

    // always @(posedge clk) begin
    //     twiddle_fac_R_add <= rom_real_data[addr];
    //     twiddle_fac_Q_add <= rom_imag_data[addr];
    //     twiddle_fac_R_sub <= rom_real_data[addr+OFFSET];
    //     twiddle_fac_Q_sub <= rom_imag_data[addr+OFFSET];
    // end

    assign twiddle_fac_R_add = rom_real_data[addr];
    assign twiddle_fac_Q_add = rom_imag_data[addr];
    assign twiddle_fac_R_sub = rom_real_data[addr+OFFSET];
    assign twiddle_fac_Q_sub = rom_imag_data[addr+OFFSET];

endmodule
